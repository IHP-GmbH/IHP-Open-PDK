************************************************************************
*
* Copyright 2024 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL sub!:G

*.PIN sub!

************************************************************************
* Library Name: sg13g2_iocell
* Cell Type:    Fillers
************************************************************************

* sg13g2_Corner
.SUBCKT sg13g2_Corner vss vdd iovss iovdd

.ENDS

* sg13g2_Filler400
.SUBCKT sg13g2_Filler400 vss vdd iovss iovdd

.ENDS

* sg13g2_Filler1000
.SUBCKT sg13g2_Filler1000 vss vdd iovss iovdd

.ENDS

* sg13g2_Filler2000
.SUBCKT sg13g2_Filler2000 vss vdd iovss iovdd

.ENDS

* sg13g2_Filler4000
.SUBCKT sg13g2_Filler4000 vss vdd iovss iovdd

.ENDS

* sg13g2_Filler10000
.SUBCKT sg13g2_Filler10000 vss vdd iovss iovdd

.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_SecondaryProtection
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_SecondaryProtection core minus pad plus
RR0 pad core 586.899 $SUB=sub! $[res_rppd] m=1 l=2u w=1u ps=180n trise=0.0 b=0
DD0 sub! core dantenna m=1 w=780n l=3.1u a=2.418p p=7.76u
XR1 minus sub! / ptap1 r=46.556 A=9.03p Perim=12.02u w=3.005u l=3.005u
DD1 core plus dpantenna m=1 w=780.00n l=4.98u a=3.884p p=11.52u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_Clamp_N20N0D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N20N0D iovss pad
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=88.000u l=600.0n ng=20
XR0 iovss sub! / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
RR1 iovss net2 1.959K $SUB=sub! $[res_rppd] m=1 l=3.54u w=500n ps=180n 
+ trise=0.0 b=0
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_Clamp_P20N0D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P20N0D iovdd iovss pad
MP0 pad net2 iovdd iovdd sg13_hv_pmos m=1 w=266.4u l=600.0n ng=40
RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
XR1 iovss sub! / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_DCNDiode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_DCNDiode anode cathode guard
DD0 sub! cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 anode sub! / ptap1 r=6.374 A=111.514p Perim=42.24u w=10.56u l=10.56u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_DCPDiode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_DCPDiode anode cathode guard
DD0 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 guard sub! / ptap1 r=17.289 A=33.524p Perim=23.16u w=5.79u l=5.79u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadAnalog
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadAnalog iovdd iovss pad padres vdd vss
XI6 padres iovss pad iovdd / sg13g2_SecondaryProtection
XI8 iovss pad / sg13g2_Clamp_N20N0D
XI9 iovdd iovss pad / sg13g2_Clamp_P20N0D
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=22.579 A=23.863p Perim=19.54u w=4.885u l=4.885u
XR2 iovss sub! / ptap1 r=214.8m A=4.3n Perim=262.3u w=65.575u l=65.575u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_LevelDown
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelDown core iovdd iovss pad vdd vss
MP0 net2 net4 vdd vdd sg13_hv_pmos m=1 w=4.65u l=450.00n ng=1
MN0 net2 net4 vss sub! sg13_hv_nmos m=1 w=2.65u l=450.00n ng=1
MN1 core net2 vss sub! sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP1 core net2 vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
XR0 vss sub! / ptap1 r=127.332 A=2.016p Perim=5.68u w=1.42u l=1.42u
XI0 net4 iovss pad iovdd / sg13g2_SecondaryProtection
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadIn
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIn iovdd iovss p2c pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI1 p2c iovdd iovss pad vdd vss / sg13g2_LevelDown
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=26.653 A=19.228p Perim=17.54u w=4.385u l=4.385u
XR2 iovss sub! / ptap1 r=173.674m A=5.35n Perim=292.58u w=73.145u l=73.145u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_io_nand2_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_nand2_x1 i0 i1 nq vdd vss
MP1 nq i1 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MP0 nq i0 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MN1 net1 i0 vss sub! sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MN0 nq i1 net1 sub! sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
XR0 vss sub! / ptap1 r=262.847 A=608.4f Perim=3.12u w=780.00n l=780.00n
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_io_inv_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_inv_x1 i nq vdd vss
MN0 nq i vss sub! sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MP0 nq i vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
XR0 vss sub! / ptap1 r=262.847 A=608.4f Perim=3.12u w=780n l=780n
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_LevelUp
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelUp i iovdd o vdd vss
MN0 net2 i vss sub! sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP0 net2 i vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
MN3 o net4 vss sub! sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN2 net4 i vss sub! sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN1 net3 net2 vss sub! sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MP3 o net4 iovdd iovdd sg13_hv_pmos m=1 w=3.9u l=450.00n ng=1
MP2 net3 net4 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
MP1 net4 net3 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
XR1 vss sub! / ptap1 r=207.099 A=912.025f Perim=3.82u w=955n l=955n
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_io_tie
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_tie vdd vss
XR0 vss sub! / ptap1 r=262.847 A=608.4f Perim=3.12u w=780.00n l=780.00n
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_io_nor2_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_nor2_x1 i0 i1 nq vdd vss
MN0 nq i0 vss sub! sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MN1 nq i1 vss sub! sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MP1 net1 i0 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MP0 nq i1 net1 vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
XR0 vss sub! / ptap1 r=262.847 A=608.4f Perim=3.12u w=780.00n l=780.00n
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_GateDecode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_GateDecode core en iovdd ngate pgate vdd vss
XI1 core en net2 vdd vss / sg13g2_io_nand2_x1
XI2 en net3 vdd vss / sg13g2_io_inv_x1
XI4 net4 iovdd ngate vdd vss / sg13g2_LevelUp
XI3 net2 iovdd pgate vdd vss / sg13g2_LevelUp
XI5 vdd vss / sg13g2_io_tie
XI0 core net3 net4 vdd vss / sg13g2_io_nor2_x1
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadInOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut30mA c2p c2p_en iovdd iovss p2c pad vdd vss
XI1 p2c iovdd iovss pad vdd vss / sg13g2_LevelDown
XI3 iovss pad iovdd / sg13g2_DCNDiode
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=66.000u l=600.0n ng=15
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=199.8u l=600.0n ng=30
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=50.701 A=8.009p Perim=11.32u w=2.83u l=2.83u
XR2 iovss sub! / ptap1 r=209.125m A=4.42n Perim=265.94u w=66.485u l=66.485u
XI0 c2p c2p_en iovdd net2 net1 vdd vss / sg13g2_GateDecode
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadInOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut4mA c2p c2p_en iovdd iovss p2c pad vdd vss
XI1 p2c iovdd iovss pad vdd vss / sg13g2_LevelDown
XI3 iovss pad iovdd / sg13g2_DCNDiode
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=8.8u l=600.0n ng=2
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=26.64u l=600.0n ng=4
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=52.392 A=7.645p Perim=11.06u w=2.765u l=2.765u
XR0 iovss sub! / ptap1 r=209.125m A=4.42n Perim=265.94u w=66.485u l=66.485u
XI0 c2p c2p_en iovdd net2 net1 vdd vss / sg13g2_GateDecode
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadInOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut16mA c2p c2p_en iovdd iovss p2c pad vdd vss
XI1 p2c iovdd iovss pad vdd vss / sg13g2_LevelDown
XI3 iovss pad iovdd / sg13g2_DCNDiode
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=35.2u l=600.0n ng=8
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=106.56u l=600.0n ng=16
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=47.799 A=8.703p Perim=11.8u w=2.95u l=2.95u
XR0 iovss sub! / ptap1 r=207.756m A=4.45n Perim=266.84u w=66.71u l=66.71u
XI0 c2p c2p_en iovdd net2 net1 vdd vss / sg13g2_GateDecode
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_LevelUpInv
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelUpInv i iovdd o vdd vss
MN0 net2 i vss sub! sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP0 net2 i vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
MN3 o net4 vss sub! sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN2 net4 net2 vss sub! sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN1 net3 i vss sub! sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MP3 o net4 iovdd iovdd sg13_hv_pmos m=1 w=3.9u l=450.00n ng=1
MP2 net3 net4 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
MP1 net4 net3 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
XR0 vss sub! / ptap1 r=190.268 A=1.051p Perim=4.1u w=1.025u l=1.025u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_GateLevelUpInv
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_GateLevelUpInv core iovdd ngate pgate vdd vss
XI1 core iovdd pgate vdd vss / sg13g2_LevelUpInv
XI0 core iovdd ngate vdd vss / sg13g2_LevelUpInv
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut16mA c2p iovdd iovss pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI6 c2p iovdd net2 net1 vdd vss / sg13g2_GateLevelUpInv
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=35.2u l=600.0n ng=8
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=106.56u l=600.0n ng=16
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=25.665 A=20.205p Perim=17.98u w=4.495u l=4.495u
XR2 iovss sub! / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut30mA c2p iovdd iovss pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI6 c2p iovdd net2 net1 vdd vss / sg13g2_GateLevelUpInv
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=66.000u l=600.0n ng=15
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=199.8u l=600.0n ng=30
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=25.534 A=20.34p Perim=18.04u w=4.51u l=4.51u
XR2 iovss sub! / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadTriOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut4mA c2p c2p_en iovdd iovss pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI7 c2p c2p_en iovdd net2 net1 vdd vss / sg13g2_GateDecode
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=8.8u l=600.0n ng=2
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=26.64u l=600.0n ng=4
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=26.152 A=19.714p Perim=17.76u w=4.44u l=4.44u
XR2 iovss sub! / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadTriOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut30mA c2p c2p_en iovdd iovss pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI7 c2p c2p_en iovdd net2 net1 vdd vss / sg13g2_GateDecode
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=66.000u l=600.0n ng=15
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=199.8u l=600.0n ng=30
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=26.561 A=19.316p Perim=17.58u w=4.395u l=4.395u
XR2 iovss sub! / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadTriOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut16mA c2p c2p_en iovdd iovss pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI7 c2p c2p_en iovdd net2 net1 vdd vss / sg13g2_GateDecode
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=35.2u l=600.0n ng=8
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=106.56u l=600.0n ng=16
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=25.84 A=20.026p Perim=17.9u w=4.475u l=4.475u
XR2 iovss sub! / ptap1 r=208.211m A=4.44n Perim=266.54u w=66.635u l=66.635u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut4mA c2p iovdd iovss pad vdd vss
XI3 iovss pad iovdd / sg13g2_DCNDiode
XI6 c2p iovdd net2 net1 vdd vss / sg13g2_GateLevelUpInv
MN0 pad net2 iovss sub! sg13_hv_nmos m=1 w=8.8u l=600.0n ng=2
MP0 pad net1 iovdd iovdd sg13_hv_pmos m=1 w=26.64u l=600.0n ng=4
XI2 pad iovdd iovss / sg13g2_DCPDiode
XR1 vss sub! / ptap1 r=26.7 A=19.184p Perim=17.52u w=4.38u l=4.38u
XR2 iovss sub! / ptap1 r=207.756m A=4.45n Perim=266.84u w=66.71u l=66.71u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_RCClampInverter
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_RCClampInverter in iovss out supply
MN1 iovss in iovss sub! sg13_hv_nmos m=1 w=126.000u l=9.5u ng=14
MN0 out in iovss sub! sg13_hv_nmos m=1 w=108.000u l=500.0n ng=12
XR0 iovss sub! / ptap1 r=9.59 A=68.973p Perim=33.22u w=8.305u l=8.305u
MP0 out in supply supply sg13_hv_pmos m=1 w=350.000u l=500.0n ng=50
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_RCClampResistor
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_RCClampResistor pin1 pin2
RR29 net15 net16 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR28 net20 net21 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR27 net23 net24 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR26 net26 net27 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR25 net29 pin2 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR24 net17 net18 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR23 net16 net17 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR22 net28 net29 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR21 net25 net26 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR20 net22 net23 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR19 net19 net20 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR18 net27 net28 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR17 net24 net25 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR16 net21 net22 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR15 net18 net19 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR14 net5 net6 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR13 net8 net9 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR12 net11 net12 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR11 net14 net15 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR10 net2 net3 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR9 net1 net2 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR8 net13 net14 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR7 net10 net11 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR6 net7 net8 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR5 net4 net5 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR4 net12 net13 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR3 net9 net10 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR2 net6 net7 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR1 net3 net4 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR0 pin1 net1 5.239K $SUB=sub! $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_Clamp_N43N43D4R
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N43N43D4R gate pad sg13g2_io_tie
MN0<1> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<2> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<3> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<4> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<5> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<6> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<7> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<8> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<9> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<10> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<11> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<12> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<13> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<14> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<15> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<16> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<17> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<18> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<19> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<20> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<21> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<22> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<23> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<24> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<25> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<26> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<27> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<28> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<29> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<30> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<31> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<32> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<33> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<34> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<35> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<36> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<37> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<38> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<39> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<40> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<41> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<42> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<43> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<44> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<45> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<46> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<47> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<48> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<49> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<50> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<51> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<52> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<53> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<54> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<55> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<56> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<57> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<58> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<59> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<60> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<61> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<62> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<63> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<64> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<65> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<66> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<67> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<68> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<69> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<70> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<71> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<72> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<73> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<74> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<75> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<76> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<77> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<78> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<79> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<80> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<81> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<82> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<83> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<84> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<85> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<86> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<87> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<88> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<89> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<90> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<91> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<92> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<93> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<94> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<95> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<96> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<97> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<98> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<99> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<100> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<101> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<102> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<103> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<104> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<105> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<106> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<107> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<108> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<109> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<110> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<111> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<112> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<113> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<114> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<115> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<116> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<117> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<118> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<119> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<120> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<121> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<122> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<123> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<124> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<125> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<126> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<127> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<128> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<129> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<130> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<131> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<132> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<133> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<134> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<135> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<136> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<137> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<138> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<139> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<140> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<141> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<142> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<143> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<144> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<145> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<146> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<147> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<148> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<149> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<150> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<151> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<152> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<153> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<154> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<155> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<156> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<157> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<158> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<159> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<160> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<161> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<162> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<163> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<164> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<165> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<166> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<167> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<168> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<169> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<170> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<171> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<172> pad gate sg13g2_io_tie sub! sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
XR0 sg13g2_io_tie sub! / ptap1 r=439m A=2.051n Perim=181.16u w=45.29u l=45.29u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadIOVdd
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIOVdd iovdd iovss vdd vss
XI1 net1 iovss net2 iovdd / sg13g2_RCClampInverter
XI2 iovdd net1 / sg13g2_RCClampResistor
XR0 vss sub! / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
XI0 net2 iovdd iovss / sg13g2_Clamp_N43N43D4R
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadIOVss
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIOVss iovdd iovss vdd vss
DD2 sub! iovss dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD1 iovss iovdd dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR2 vss sub! / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XR0 iovss sub! / ptap1 r=169.45m A=5.487n Perim=296.3u w=74.075u l=74.075u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadVdd
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadVdd iovdd iovss vdd vss
DD1 vdd iovdd dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 vss sub! / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XR1 iovss sub! / ptap1 r=168.319m A=5.525n Perim=297.32u w=74.33u l=74.33u
DD0 sub! vdd dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
.ENDS

************************************************************************
* Library Name: sg13g2_iocell
* Cell Name:    sg13g2_IOPadVss
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadVss iovdd iovss vdd vss
XI1 iovss vss iovss / sg13g2_DCNDiode
XI2 vss iovdd iovss / sg13g2_DCPDiode
XR1 iovss sub! / ptap1 r=174.346m A=5.329n Perim=292u w=73u l=73u
XR0 vss sub! / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS


