************************************************************************
* 
* Copyright 2023 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
************************************************************************

.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_CORNER VDD_CORE VSS
XI16 VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR LWL NW PW VDD VSS
MN1 VSS LWL VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 VSS net9 VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR A_WL<15> A_WL<14> A_WL<13> A_WL<12> 
+ A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> 
+ A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS
XI0<15> A_WL<15> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<14> A_WL<14> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<13> A_WL<13> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<12> A_WL<12> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<11> A_WL<11> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<10> A_WL<10> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<9> A_WL<9> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<8> A_WL<8> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<7> A_WL<7> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<6> A_WL<6> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<5> A_WL<5> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<4> A_WL<4> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<3> A_WL<3> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<2> A_WL<2> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<1> A_WL<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
XI0<0> A_WL<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_LR
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL BLC_BOT BLC_TOP BLT_BOT BLT_TOP LWL NW PW 
+ RWL VDD VSS
MN0 NC NT VSS PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN1 NT NC VSS PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN3 NC RWL BLC_TOP PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN2 BLT_BOT LWL NT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 NT NC VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 NC NT VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
R1 BLC_BOT BLC_TOP lvsres w=2.6e-07 l=6e-07
R0 BLT_BOT BLT_TOP lvsres w=2.6e-07 l=6e-07
R2 RWL LWL lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> 
+ A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<15> 
+ A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> 
+ A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> 
+ A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> 
+ A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE 
+ VSS
XCELL<31> A_BLC_TOP<1> A_RBLC<15> A_BLT_TOP<1> A_RBLT<15> A_RWL<15> 
+ VDD_CORE VSS A_XWL<15> VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<30> A_RBLC<14> A_RBLC<15> A_RBLT<14> A_RBLT<15> A_RWL<14> VDD_CORE 
+ VSS A_XWL<14> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<29> A_RBLC<14> A_RBLC<13> A_RBLT<14> A_RBLT<13> A_RWL<13> VDD_CORE 
+ VSS A_XWL<13> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<28> A_RBLC<12> A_RBLC<13> A_RBLT<12> A_RBLT<13> A_RWL<12> VDD_CORE 
+ VSS A_XWL<12> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<27> A_RBLC<12> A_RBLC<11> A_RBLT<12> A_RBLT<11> A_RWL<11> VDD_CORE 
+ VSS A_XWL<11> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<26> A_RBLC<10> A_RBLC<11> A_RBLT<10> A_RBLT<11> A_RWL<10> VDD_CORE 
+ VSS A_XWL<10> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<25> A_RBLC<10> A_RBLC<9> A_RBLT<10> A_RBLT<9> A_RWL<9> VDD_CORE 
+ VSS A_XWL<9> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<24> A_RBLC<8> A_RBLC<9> A_RBLT<8> A_RBLT<9> A_RWL<8> VDD_CORE 
+ VSS A_XWL<8> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<23> A_RBLC<8> A_RBLC<7> A_RBLT<8> A_RBLT<7> A_RWL<7> VDD_CORE 
+ VSS A_XWL<7> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<22> A_RBLC<6> A_RBLC<7> A_RBLT<6> A_RBLT<7> A_RWL<6> VDD_CORE 
+ VSS A_XWL<6> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<21> A_RBLC<6> A_RBLC<5> A_RBLT<6> A_RBLT<5> A_RWL<5> VDD_CORE 
+ VSS A_XWL<5> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<20> A_RBLC<4> A_RBLC<5> A_RBLT<4> A_RBLT<5> A_RWL<4> VDD_CORE 
+ VSS A_XWL<4> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<19> A_RBLC<4> A_RBLC<3> A_RBLT<4> A_RBLT<3> A_RWL<3> VDD_CORE 
+ VSS A_XWL<3> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<18> A_RBLC<2> A_RBLC<3> A_RBLT<2> A_RBLT<3> A_RWL<2> VDD_CORE 
+ VSS A_XWL<2> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<17> A_RBLC<2> A_RBLC<1> A_RBLT<2> A_RBLT<1> A_RWL<1> VDD_CORE 
+ VSS A_XWL<1> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<16> A_BLC_BOT<1> A_RBLC<1> A_BLT_BOT<1> A_RBLT<1> A_RWL<0> VDD_CORE 
+ VSS A_XWL<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<15> A_BLC_TOP<0> A_LBLC<15> A_BLT_TOP<0> A_LBLT<15> A_LWL<15> 
+ VDD_CORE VSS A_XWL<15> VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<14> A_LBLC<14> A_LBLC<15> A_LBLT<14> A_LBLT<15> A_LWL<14> VDD_CORE 
+ VSS A_XWL<14> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<13> A_LBLC<14> A_LBLC<13> A_LBLT<14> A_LBLT<13> A_LWL<13> VDD_CORE 
+ VSS A_XWL<13> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<12> A_LBLC<12> A_LBLC<13> A_LBLT<12> A_LBLT<13> A_LWL<12> VDD_CORE 
+ VSS A_XWL<12> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<11> A_LBLC<12> A_LBLC<11> A_LBLT<12> A_LBLT<11> A_LWL<11> VDD_CORE 
+ VSS A_XWL<11> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<10> A_LBLC<10> A_LBLC<11> A_LBLT<10> A_LBLT<11> A_LWL<10> VDD_CORE 
+ VSS A_XWL<10> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<9> A_LBLC<10> A_LBLC<9> A_LBLT<10> A_LBLT<9> A_LWL<9> VDD_CORE 
+ VSS A_XWL<9> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<8> A_LBLC<8> A_LBLC<9> A_LBLT<8> A_LBLT<9> A_LWL<8> VDD_CORE 
+ VSS A_XWL<8> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<7> A_LBLC<8> A_LBLC<7> A_LBLT<8> A_LBLT<7> A_LWL<7> VDD_CORE 
+ VSS A_XWL<7> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<6> A_LBLC<6> A_LBLC<7> A_LBLT<6> A_LBLT<7> A_LWL<6> VDD_CORE 
+ VSS A_XWL<6> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<5> A_LBLC<6> A_LBLC<5> A_LBLT<6> A_LBLT<5> A_LWL<5> VDD_CORE 
+ VSS A_XWL<5> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<4> A_LBLC<4> A_LBLC<5> A_LBLT<4> A_LBLT<5> A_LWL<4> VDD_CORE 
+ VSS A_XWL<4> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<3> A_LBLC<4> A_LBLC<3> A_LBLT<4> A_LBLT<3> A_LWL<3> VDD_CORE 
+ VSS A_XWL<3> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<2> A_LBLC<2> A_LBLC<3> A_LBLT<2> A_LBLT<3> A_LWL<2> VDD_CORE 
+ VSS A_XWL<2> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<1> A_LBLC<2> A_LBLC<1> A_LBLT<2> A_LBLT<1> A_LWL<1> VDD_CORE 
+ VSS A_XWL<1> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
XCELL<0> A_BLC_BOT<0> A_LBLC<1> A_BLT_BOT<0> A_LBLT<1> A_LWL<0> VDD_CORE 
+ VSS A_XWL<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_CELL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB BLC BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_TB A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ VDD_CORE VSS
XEDGE<1> A_BLC<1> A_BLT<1> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB
XEDGE<0> A_BLC<0> A_BLT<0> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB
.ENDS

.SUBCKT RSC_IHPSG13_CBUFX4 A Z VDD VSS
MN0 net9 A VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 Z net9 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP0 net9 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 Z net9 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDRV13X4 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX4 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net6 A VSS VSS nmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_WLDRV16X4 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX4
.ENDS
.SUBCKT RSC_IHPSG13_FILLCAP8 VDD VSS
MN0 vss_r vdd_r VSS VSS nmos m=1 w=4.98u l=130.00n ng=6 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD pmos m=1 w=6.48u l=385.000n ng=4 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_LHPQX2 CP D Q VDD VSS
MN3 QIN CPN net14 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN2 net14 net10 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN5 net21 D VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 QIN CP net21 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net10 QIN VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 CPN CP VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 Q QIN VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP2 QIN CP net16 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 CPN CP VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 Q QIN VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP3 net10 QIN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net16 net10 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP6 QIN CPN net20 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP5 net20 D VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NAND2X2 A B Z VDD VSS
MP1 Z B VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN0 Z B net7 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net7 A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX4 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX2 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_INVX2 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NAND3X2 A B C Z VDD VSS
MP2 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 Z B VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z C VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN1 net12 B net16 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN0 Z C net12 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN2 net16 A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NOR3X2 A B C Z VDD VSS
MP0 net13 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP2 Z C net10 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 net10 B net13 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN1 Z B VSS VSS nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
MN0 Z C VSS VSS nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
MN2 Z A VSS VSS nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_FILLCAP4 VDD VSS
MN0 vss_r vdd_r VSS VSS nmos m=1 w=2.49u l=130.00n ng=3 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD pmos m=1 w=3.24u l=385.000n ng=2 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MET2RES A B
R0 B A lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_DEC04 ADDR<3> ADDR<2> ADDR<1> ADDR<0> CS ECLK_H_BOT 
+ ECLK_H_TOP ECLK_L_BOT ECLK_L_TOP WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> 
+ WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> VDD VSS
XLATCH<3> CS ADDR<3> PADR<3> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<2> CS ADDR<2> PADR<2> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<1> CS ADDR<1> PADR<1> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<0> CS ADDR<0> PADR<0> VDD VSS / RSC_IHPSG13_LHPQX2
XI0<3> PADR<1> PADR<0> sel01<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<2> PADR<1> NADR<0> sel01<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<1> NADR<1> PADR<0> sel01<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<0> NADR<1> NADR<0> sel01<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI4 ECLK_L_BOT EN VDD VSS / RSC_IHPSG13_CINVX4
XI5 ECLK_H_BOT ECLK_L_BOT VDD VSS / RSC_IHPSG13_CINVX2
XI3<3> PADR<3> NADR<3> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> PADR<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> PADR<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> PADR<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1<3> PADR<2> PADR<3> CS sel23<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<2> PADR<3> CS sel23<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<2> NADR<3> CS sel23<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<2> NADR<3> CS sel23<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI2<15> sel23<3> sel01<3> EN WL<15> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<14> sel23<3> sel01<2> EN WL<14> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<13> sel23<3> sel01<1> EN WL<13> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<12> sel23<3> sel01<0> EN WL<12> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<11> sel23<2> sel01<3> EN WL<11> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<10> sel23<2> sel01<2> EN WL<10> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<9> sel23<2> sel01<1> EN WL<9> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<8> sel23<2> sel01<0> EN WL<8> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<7> sel23<1> sel01<3> EN WL<7> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<6> sel23<1> sel01<2> EN WL<6> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<5> sel23<1> sel01<1> EN WL<5> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<4> sel23<1> sel01<0> EN WL<4> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<3> sel23<0> sel01<3> EN WL<3> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<2> sel23<0> sel01<2> EN WL<2> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<1> sel23<0> sel01<1> EN WL<1> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<0> sel23<0> sel01<0> EN WL<0> VDD VSS / RSC_IHPSG13_NOR3X2
XCAPS4 VDD VSS / RSC_IHPSG13_FILLCAP4
XI11 ECLK_L_BOT ECLK_L_TOP / RSC_IHPSG13_MET2RES
XR0 ECLK_H_BOT ECLK_H_TOP / RSC_IHPSG13_MET2RES
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWDEC4 ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> 
+ CS_I ECLK_I WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XSEL ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I ECLK_H<1> 
+ ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> 
+ WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> 
+ WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
.ENDS
.SUBCKT RSC_IHPSG13_CINVX8 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=2.82u l=130.00n ng=4 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_DFNQMX2IX1 BE BI CN D QI QIN VDD VSS
MN15 net026 BI VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN14 MXI_OUT BE net026 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net025 D VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 MXI_OUT BEN net025 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN10 QI CNN net21 VSS nmos m=1 w=850.00n l=130.00n ng=1 nrd=0 nrs=0
MN11 net21 QI_MS VSS VSS nmos m=1 w=850.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN7 net30 QI_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN6 QIN_MS CNN net30 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 QI_MS QIN_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN12 CNN CN VSS VSS nmos m=1 w=495.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN9 net37 MXI_OUT VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN8 QIN_MS CN net37 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 QI CN net25 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN4 net25 QIN VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 QIN QI VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN13 BEN BE VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP15 MXI_OUT BEN net027 VDD pmos m=1 w=985.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP14 net027 BI VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP1 MXI_OUT BE net024 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net024 D VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP13 BEN BE VDD VDD pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 QI_MS QIN_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP3 QI CNN net27 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MP2 net27 QIN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP10 net36 MXI_OUT VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP11 QIN_MS CNN net36 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net32 QI_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 QIN_MS CN net32 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 QIN QI VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP12 CNN CN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP9 QI CN net19 VDD pmos m=1 w=990.00n l=130.00n ng=1 nrd=0 nrs=0
MP8 net19 QI_MS VDD VDD pmos m=1 w=990.00n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWREG4 ACLK_N_I ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX1 A Z VDD VSS
MN1 net010 net032 VSS VSS nmos m=1 w=300.0n l=160.00n ng=1 
+ nrd=0 nrs=0
MN2 net032 A net014 VSS nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MN0 Z net032 net010 VSS nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MN3 net014 A VSS VSS nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MP1 Z net032 net07 VDD pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
MP3 net011 A VDD VDD pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
MP0 net07 net032 VDD VDD pmos m=1 w=720.00n l=160.00n ng=1 
+ nrd=0 nrs=0
MP2 net032 A net011 VDD pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX1_DUMMY A Z VDD VSS
MN0 vss_r vdd_r VSS VSS nmos m=1 w=2.49u l=300.0n ng=3 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD pmos m=1 w=3.24u l=640.00n ng=2 nrd=0 
+ nrs=0
R0 Z A lvsres w=2.6e-07 l=6e-07
.ENDS

.SUBCKT RSC_IHPSG13_MX2IX1 A0 A1 S ZN VDD VSS
MP4 SN S VDD VDD pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 nrs=0
MP3 ZN SN net12 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 nrs=0
MP2 net12 A1 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 ZN S net17 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 net17 A0 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 SN S VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN3 net13 A1 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 ZN S net13 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net15 A0 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 ZN SN net15 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_DLY_MUX A SEL Z VDD VSS
XI11 net4 Z VDD VSS / RSC_IHPSG13_CINVX2
XI8 A D<3> SEL net4 VDD VSS / RSC_IHPSG13_MX2IX1
XI20<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1
.ENDS
.SUBCKT RSC_IHPSG13_DFNQX2 CN D Q VDD VSS
MN0 Q QIN_SL VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN10 QIN_SL CNN net21 VSS nmos m=1 w=850.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN11 net21 QI_MS VSS VSS nmos m=1 w=850.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN7 net30 QI_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN6 QIN_MS CNN net30 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 QI_MS QIN_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN12 CNN CN VSS VSS nmos m=1 w=495.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN9 net37 D VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN8 QIN_MS CN net37 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 QIN_SL CN net25 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net25 QI_SL VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN2 QI_SL QIN_SL VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP0 Q QIN_SL VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 QI_MS QIN_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP3 QIN_SL CNN net27 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net27 QI_SL VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP10 net36 D VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP11 QIN_MS CNN net36 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net32 QI_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 QIN_MS CN net32 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 QI_SL QIN_SL VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP12 CNN CN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP9 QIN_SL CN net19 VDD pmos m=1 w=990.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP8 net19 QI_MS VDD VDD pmos m=1 w=990.00n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CNAND2X2 A B Z VDD VSS
MN0 Z B net6 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net6 A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 Z B VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CGATEPX4 CP E Q VDD VSS
MN1 net08 QIN VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net019 net08 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN3 QIN CP net019 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN6 Q net015 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 
+ nrs=0
MN5 net015 net08 net018 VSS nmos m=1 w=980.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN8 QIN CPN net023 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN7 net023 E VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net018 CP VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 CPN CP VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP3 net08 QIN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 QIN CPN net017 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net017 net08 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP0 CPN CP VDD VDD pmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP8 QIN CP net024 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 net024 E VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net015 CP VDD VDD pmos m=1 w=1.27u l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 Q net015 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 
+ nrs=0
MP5 net015 net08 VDD VDD pmos m=1 w=1.27u l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CBUFX8 A Z VDD VSS
MP0 net4 A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net4 VDD VDD pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
MN1 Z net4 VSS VSS nmos m=1 w=2.82u l=130.00n ng=4 nrd=0 nrs=0
MN0 net4 A VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX2 A Z VDD VSS
MN2 net4 A net9 VSS nmos m=1 w=320.00n l=200.0n ng=1 nrd=0 nrs=0
MN0 Z net4 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net9 A VSS VSS nmos m=1 w=320.00n l=200.0n ng=1 nrd=0 nrs=0
MP2 net4 A net10 VDD pmos m=1 w=1.2u l=200.0n ng=1 nrd=0 nrs=0
MP1 net10 A VDD VDD pmos m=1 w=1.2u l=200.0n ng=1 nrd=0 nrs=0
MP0 Z net4 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MX2X2 A0 A1 S Z VDD VSS
MP6 Z net010 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 SN S VDD VDD pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 nrs=0
MP3 net010 SN net12 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net12 A1 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net010 S net17 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net17 A0 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 Z net010 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 SN S VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 nrs=0
MN3 net13 A1 VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net010 S net13 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net15 A0 VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net010 SN net15 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_AND2X2 A B Z VDD VSS
MN3 Z net6 VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net9 B VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net6 B VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_TIEL Z VDD VSS
MN0 Z net2 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net2 net2 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_XOR2X2 A B Z VDD VSS
MP8 net012 B net7 VDD pmos m=1 w=825.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 net011 net3 net012 VDD pmos m=1 w=825.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP6 Z net012 VDD VDD pmos m=1 w=1.535u l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net7 A VDD VDD pmos m=1 w=825.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net011 net7 VDD VDD pmos m=1 w=825.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 net3 B VDD VDD pmos m=1 w=580.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN7 net012 B net011 VSS nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 net7 net3 net012 VSS nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 Z net012 VSS VSS nmos m=1 w=775.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net7 A VSS VSS nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net3 B VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 net011 net7 VSS VSS nmos m=1 w=555.000n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_OA12X1 A B C Z VDD VSS
MN2 net7 C VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 Z net17 VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net17 B net7 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN0 net17 A net7 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 net24 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP3 Z net17 VDD VDD pmos m=1 w=905.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net17 B net24 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP2 net17 C VDD VDD pmos m=1 w=905.000n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_CTRL ACLK_N BIST_CK_I BIST_CS_I BIST_EN BIST_RE_I 
+ BIST_WE_I B_TIEL_O CK_I CS_I DCLK ECLK PULSE_H PULSE_L PULSE_O RCLK RE_I 
+ ROW_CS WCLK WE_I VDD VSS
XI17 ck_regs we col_we VDD VSS / RSC_IHPSG13_DFNQX2
XI16 ck_regs re col_re VDD VSS / RSC_IHPSG13_DFNQX2
XI18 ck_regs cs net7 VDD VSS / RSC_IHPSG13_DFNQX2
XI71 ACLK_N net012 PULSE_O VDD VSS / RSC_IHPSG13_DFNQX2
XI77 col_we net9 net016 VDD VSS / RSC_IHPSG13_CNAND2X2
XI76 col_re net9 net018 VDD VSS / RSC_IHPSG13_CNAND2X2
XI15 ck_dly WEorREandCS aclk VDD VSS / RSC_IHPSG13_CGATEPX4
XI14 ck WEandCS DCLK VDD VSS / RSC_IHPSG13_CGATEPX4
XI60 net7 ROW_CS VDD VSS / RSC_IHPSG13_CBUFX8
XI73 PULSE_O net012 VDD VSS / RSC_IHPSG13_CINVX2
XI8 net9 net8 VDD VSS / RSC_IHPSG13_CINVX2
XI64 ck ck_dly VDD VSS / RSC_IHPSG13_CDLYX2
XI86 CS_I BIST_CS_I BIST_EN cs VDD VSS / RSC_IHPSG13_MX2X2
XI87 CK_I BIST_CK_I BIST_EN ck VDD VSS / RSC_IHPSG13_MX2X2
XI85 WE_I BIST_WE_I BIST_EN we VDD VSS / RSC_IHPSG13_MX2X2
XI84 RE_I BIST_RE_I BIST_EN re VDD VSS / RSC_IHPSG13_MX2X2
XI22 we cs WEandCS VDD VSS / RSC_IHPSG13_AND2X2
XBM_TIEL B_TIEL_O VDD VSS / RSC_IHPSG13_TIEL
XI48 ck_dly ck_regs VDD VSS / RSC_IHPSG13_CINVX4
XI81 net016 WCLK VDD VSS / RSC_IHPSG13_CINVX4
XI80 net018 RCLK VDD VSS / RSC_IHPSG13_CINVX4
XI78 net8 net020 VDD VSS / RSC_IHPSG13_CINVX4
XI6 PULSE_L PULSE_H net9 VDD VSS / RSC_IHPSG13_XOR2X2
XI79 net020 ECLK VDD VSS / RSC_IHPSG13_CINVX8
XI63 aclk ACLK_N VDD VSS / RSC_IHPSG13_CINVX8
XI21 re we cs WEorREandCS VDD VSS / RSC_IHPSG13_OA12X1
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDEC2 ACLK_N ADDR<1> ADDR<0> ADDR_COL<1> ADDR_COL<0> 
+ ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> ADDR_DEC<2> 
+ ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI14<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net6<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net6<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<3> PADR<1> PADR<0> addr_n<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<2> PADR<1> NADR<0> addr_n<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<1> NADR<1> PADR<0> addr_n<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<0> NADR<1> NADR<0> addr_n<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI16<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI17<3> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_TIEL
XI17<2> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_TIEL
XI17<1> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_TIEL
XI17<0> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RSC_IHPSG13_NOR2X2 A B Z VDD VSS
MP1 Z B net9 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net9 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN0 Z B VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 Z A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX4_WN A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BLDRV BLC BLC_SEL BLT BLT_SEL PRE_N SEL_P WR_ONE WR_ZERO 
+ VDD VSS
XCDEC SEL_P WR_ZERO BLC_PMOS_DRIVE VDD VSS / RSC_IHPSG13_NAND2X2
XTDEC SEL_P WR_ONE BLT_PMOS_DRIVE VDD VSS / RSC_IHPSG13_NAND2X2
MTWN BLT BLT_NMOS_DRIVE VSS VSS nmos m=1 w=4.82u l=130.00n 
+ ng=2 nrd=0 nrs=0
MCWN BLC BLC_NMOS_DRIVE VSS VSS nmos m=1 w=4.82u l=130.00n 
+ ng=2 nrd=0 nrs=0
MCWP BLC BLC_PMOS_DRIVE VDD VDD pmos m=1 w=1.5u l=130.00n ng=1 
+ nrd=0 nrs=0
MTWP BLT BLT_PMOS_DRIVE VDD VDD pmos m=1 w=1.5u l=130.00n ng=1 
+ nrd=0 nrs=0
MTSP BLT_SEL SEL_N BLT VDD pmos m=1 w=1.5u l=130.00n ng=1 nrd=0 
+ nrs=0
MTPR BLT PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n ng=2 nrd=0 
+ nrs=0
MCSP BLC_SEL SEL_N BLC VDD pmos m=1 w=1.5u l=130.00n ng=1 nrd=0 
+ nrs=0
MCPR BLC PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n ng=2 nrd=0 
+ nrs=0
XI86 SEL_P SEL_N VDD VSS / RSC_IHPSG13_INVX2
XTINV BLC_PMOS_DRIVE BLT_NMOS_DRIVE VDD VSS / RSC_IHPSG13_INVX2
XCINV BLT_PMOS_DRIVE BLC_NMOS_DRIVE VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RSC_IHPSG13_TIEH Z VDD VSS
MN0 net2 net2 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 Z net2 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MET3RES A B
R0 B A lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RSC_IHPSG13_DFPQD_MSAFFX2 CP DN DP QN QP VDD VSS
MN12 SN RN DIFFP VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN13 TAIL CP VSS VSS nmos m=1 w=2.4u l=130.00n ng=2 nrd=0 nrs=0
MN9 DIFFP DP TAIL VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN10 DIFFN DN TAIL VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN11 RN SN DIFFN VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN19 net33 SN VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN20 QN QP net37 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN18 net37 RN VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN17 QP QN net33 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP15 SN RN VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP16 RN CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP14 DIFFP CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MP12 RN SN VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP13 DIFFN CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MP11 SN CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP19 QN QP VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
MP20 QP SN VDD VDD pmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP18 QN RN VDD VDD pmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP17 QP QN VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CBUFX2 A Z VDD VSS
MN1 Z net4 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net4 A VSS VSS nmos m=1 w=540.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 Z net4 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net4 A VDD VDD pmos m=1 w=1.1u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_INVX4 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=1.96u l=130.00n ng=2 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLCTRL2 A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<3> A_BLC<2> A_BLC<1> 
+ A_BLC<0> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I80 A_WCLK_B_R A_RCLK_B_R net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I44 A_WCLK_B_R A_BM_N A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_ADDR_DEC<2> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_ADDR_DEC<1> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<0> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_R A_RCLK_B_L / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_R A_RCLK_L / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_R A_WCLK_B_L / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I78 A_RCLK_B_R A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_R VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_R A_RCLK_B_R VDD VSS / RSC_IHPSG13_CINVX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4 VDD VSS
XI0<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2 VDD VSS
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDEC4 ACLK_N ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<3> BIST_ADDR<2> 
+ BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI15 ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI14 addr_int ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int net7<0> VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RSC_IHPSG13_AND2X4 A B Z VDD VSS
MN3 Z net6 VSS VSS nmos m=1 w=1.96u l=130.00n ng=2 nrd=0 nrs=0
MN4 net9 B VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP0 net6 B VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLCTRL4 A_ADDR_COL A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<15> A_BLC<14> 
+ A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> 
+ A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> 
+ A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L 
+ A_DCLK_B_R A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L 
+ A_RCLK_R A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_I80 A_WCLK_B_L A_RCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DO_WRITE_P A_DI_N A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XA_CAPS<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_N0 A_P0 VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL A_N0 VDD VSS / RSC_IHPSG13_CINVX4
XA_I81<1> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<15> A_BLC<15> A_BLC_SEL A_BLT<15> A_BLT_SEL A_PRE_N A_SEL_P<15> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<14> A_BLC<14> A_BLC_SEL A_BLT<14> A_BLT_SEL A_PRE_N A_SEL_P<14> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<13> A_BLC<13> A_BLC_SEL A_BLT<13> A_BLT_SEL A_PRE_N A_SEL_P<13> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<12> A_BLC<12> A_BLC_SEL A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<12> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<11> A_BLC<11> A_BLC_SEL A_BLT<11> A_BLT_SEL A_PRE_N A_SEL_P<11> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<10> A_BLC<10> A_BLC_SEL A_BLT<10> A_BLT_SEL A_PRE_N A_SEL_P<10> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<9> A_BLC<9> A_BLC_SEL A_BLT<9> A_BLT_SEL A_PRE_N A_SEL_P<9> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<8> A_BLC<8> A_BLC_SEL A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<8> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_SEL_P<7> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_SEL_P<6> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_SEL_P<5> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<4> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_SEL_P<3> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_SEL_P<2> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_SEL_P<1> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<0> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net24 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3INV<15> net23<0> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<1> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<2> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<3> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<4> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<5> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<6> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<7> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<8> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<9> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<10> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<11> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<12> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<13> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<14> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<15> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I70<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_DEC3<15> A_P0 A_ADDR_DEC<7> net23<0> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<14> A_P0 A_ADDR_DEC<6> net23<1> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<13> A_P0 A_ADDR_DEC<5> net23<2> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<12> A_P0 A_ADDR_DEC<4> net23<3> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<11> A_P0 A_ADDR_DEC<3> net23<4> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<10> A_P0 A_ADDR_DEC<2> net23<5> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<9> A_P0 A_ADDR_DEC<1> net23<6> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<8> A_P0 A_ADDR_DEC<0> net23<7> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<7> A_N0 A_ADDR_DEC<7> net23<8> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<6> A_N0 A_ADDR_DEC<6> net23<9> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<5> A_N0 A_ADDR_DEC<5> net23<10> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<4> A_N0 A_ADDR_DEC<4> net23<11> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<3> A_N0 A_ADDR_DEC<3> net23<12> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<2> A_N0 A_ADDR_DEC<2> net23<13> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<1> A_N0 A_ADDR_DEC<1> net23<14> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<0> A_N0 A_ADDR_DEC<0> net23<15> VDD VSS / RSC_IHPSG13_NAND2X2
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDEC3 ACLK_N ADDR<2> ADDR<1> ADDR<0> ADDR_COL<1> 
+ ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> 
+ ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> 
+ BIST_EN_I VDD VSS
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net6<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net6<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net6<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLCTRL3 A_ADDR_DEC<7> A_ADDR_DEC<6> A_ADDR_DEC<5> 
+ A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> A_ADDR_DEC<0> 
+ A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> 
+ A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R A_DCLK_L 
+ A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R A_TIEH_O 
+ A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_R A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_I70<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I44 A_BM_N A_WCLK_B_R A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_ADDR_DEC<7> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_ADDR_DEC<6> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_ADDR_DEC<5> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_ADDR_DEC<4> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_ADDR_DEC<2> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_ADDR_DEC<1> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<0> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I80 A_WCLK_B_R A_RCLK_B_R net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_16x2_CORNER VDD_CORE VSS
XI16 VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR A_WL B_WL NW PW VDD VSS
MN1 VSS A_WL VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 VSS B_WL VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_16x2_EDGE_LR A_WL<15> A_WL<14> A_WL<13> A_WL<12> 
+ A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> 
+ A_WL<2> A_WL<1> A_WL<0> B_WL<15> B_WL<14> B_WL<13> B_WL<12> B_WL<11> 
+ B_WL<10> B_WL<9> B_WL<8> B_WL<7> B_WL<6> B_WL<5> B_WL<4> B_WL<3> B_WL<2> 
+ B_WL<1> B_WL<0> VDD_CORE VSS
XI0<15> A_WL<15> B_WL<15> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<14> A_WL<14> B_WL<14> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<13> A_WL<13> B_WL<13> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<12> A_WL<12> B_WL<12> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<11> A_WL<11> B_WL<11> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<10> A_WL<10> B_WL<10> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<9> A_WL<9> B_WL<9> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<8> A_WL<8> B_WL<8> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<7> A_WL<7> B_WL<7> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<6> A_WL<6> B_WL<6> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<5> A_WL<5> B_WL<5> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<4> A_WL<4> B_WL<4> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<3> A_WL<3> B_WL<3> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<2> A_WL<2> B_WL<2> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<1> A_WL<1> B_WL<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
XI0<0> A_WL<0> B_WL<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_LR
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL A_BLC_BOT A_BLC_TOP A_BLT_BOT A_BLT_TOP 
+ A_LWL A_RWL B_BLC_BOT B_BLC_TOP B_BLT_BOT B_BLT_TOP B_LWL B_RWL NW PW VDD VSS
MN5 NC B_RWL B_BLC_BOT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN4 B_BLT_BOT B_LWL NT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 NC NT VSS PW nmos m=1 w=600.0n l=130.00n ng=2 nrd=0 nrs=0
MN1 NT NC VSS PW nmos m=1 w=600.0n l=130.00n ng=2 nrd=0 nrs=0
MN3 NC A_RWL A_BLC_TOP PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN2 A_BLT_TOP A_LWL NT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 NT NC VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 NC NT VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
R5 B_RWL B_LWL lvsres w=2.6e-07 l=6e-07
R4 B_BLC_BOT B_BLC_TOP lvsres w=2.6e-07 l=6e-07
R3 B_BLT_BOT B_BLT_TOP lvsres w=2.6e-07 l=6e-07
R1 A_BLC_BOT A_BLC_TOP lvsres w=2.6e-07 l=6e-07
R0 A_BLT_BOT A_BLT_TOP lvsres w=2.6e-07 l=6e-07
R2 A_RWL A_LWL lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_16x2_SRAM A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> 
+ A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<15> 
+ A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> 
+ A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> 
+ A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> 
+ A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> B_BLC_BOT<1> 
+ B_BLC_BOT<0> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT_BOT<1> B_BLT_BOT<0> 
+ B_BLT_TOP<1> B_BLT_TOP<0> B_LWL<15> B_LWL<14> B_LWL<13> B_LWL<12> B_LWL<11> 
+ B_LWL<10> B_LWL<9> B_LWL<8> B_LWL<7> B_LWL<6> B_LWL<5> B_LWL<4> B_LWL<3> 
+ B_LWL<2> B_LWL<1> B_LWL<0> B_RWL<15> B_RWL<14> B_RWL<13> B_RWL<12> B_RWL<11> 
+ B_RWL<10> B_RWL<9> B_RWL<8> B_RWL<7> B_RWL<6> B_RWL<5> B_RWL<4> B_RWL<3> 
+ B_RWL<2> B_RWL<1> B_RWL<0> VDD_CORE VSS
XCELL<31> A_BLC_TOP<1> A_RBLC<15> A_BLT_TOP<1> A_RBLT<15> A_XWL<15> A_RWL<15> 
+ B_BLC_TOP<1> B_RBLC<15> B_BLT_TOP<1> B_RBLT<15> B_XWL<15> B_RWL<15> 
+ VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<30> A_RBLC<14> A_RBLC<15> A_RBLT<14> A_RBLT<15> A_XWL<14> A_RWL<14> 
+ B_RBLC<14> B_RBLC<15> B_RBLT<14> B_RBLT<15> B_XWL<14> B_RWL<14> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<29> A_RBLC<14> A_RBLC<13> A_RBLT<14> A_RBLT<13> A_XWL<13> A_RWL<13> 
+ B_RBLC<14> B_RBLC<13> B_RBLT<14> B_RBLT<13> B_XWL<13> B_RWL<13> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<28> A_RBLC<12> A_RBLC<13> A_RBLT<12> A_RBLT<13> A_XWL<12> A_RWL<12> 
+ B_RBLC<12> B_RBLC<13> B_RBLT<12> B_RBLT<13> B_XWL<12> B_RWL<12> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<27> A_RBLC<12> A_RBLC<11> A_RBLT<12> A_RBLT<11> A_XWL<11> A_RWL<11> 
+ B_RBLC<12> B_RBLC<11> B_RBLT<12> B_RBLT<11> B_XWL<11> B_RWL<11> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<26> A_RBLC<10> A_RBLC<11> A_RBLT<10> A_RBLT<11> A_XWL<10> A_RWL<10> 
+ B_RBLC<10> B_RBLC<11> B_RBLT<10> B_RBLT<11> B_XWL<10> B_RWL<10> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<25> A_RBLC<10> A_RBLC<9> A_RBLT<10> A_RBLT<9> A_XWL<9> A_RWL<9> 
+ B_RBLC<10> B_RBLC<9> B_RBLT<10> B_RBLT<9> B_XWL<9> B_RWL<9> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<24> A_RBLC<8> A_RBLC<9> A_RBLT<8> A_RBLT<9> A_XWL<8> A_RWL<8> B_RBLC<8> 
+ B_RBLC<9> B_RBLT<8> B_RBLT<9> B_XWL<8> B_RWL<8> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<23> A_RBLC<8> A_RBLC<7> A_RBLT<8> A_RBLT<7> A_XWL<7> A_RWL<7> B_RBLC<8> 
+ B_RBLC<7> B_RBLT<8> B_RBLT<7> B_XWL<7> B_RWL<7> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<22> A_RBLC<6> A_RBLC<7> A_RBLT<6> A_RBLT<7> A_XWL<6> A_RWL<6> B_RBLC<6> 
+ B_RBLC<7> B_RBLT<6> B_RBLT<7> B_XWL<6> B_RWL<6> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<21> A_RBLC<6> A_RBLC<5> A_RBLT<6> A_RBLT<5> A_XWL<5> A_RWL<5> B_RBLC<6> 
+ B_RBLC<5> B_RBLT<6> B_RBLT<5> B_XWL<5> B_RWL<5> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<20> A_RBLC<4> A_RBLC<5> A_RBLT<4> A_RBLT<5> A_XWL<4> A_RWL<4> B_RBLC<4> 
+ B_RBLC<5> B_RBLT<4> B_RBLT<5> B_XWL<4> B_RWL<4> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<19> A_RBLC<4> A_RBLC<3> A_RBLT<4> A_RBLT<3> A_XWL<3> A_RWL<3> B_RBLC<4> 
+ B_RBLC<3> B_RBLT<4> B_RBLT<3> B_XWL<3> B_RWL<3> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<18> A_RBLC<2> A_RBLC<3> A_RBLT<2> A_RBLT<3> A_XWL<2> A_RWL<2> B_RBLC<2> 
+ B_RBLC<3> B_RBLT<2> B_RBLT<3> B_XWL<2> B_RWL<2> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<17> A_RBLC<2> A_RBLC<1> A_RBLT<2> A_RBLT<1> A_XWL<1> A_RWL<1> B_RBLC<2> 
+ B_RBLC<1> B_RBLT<2> B_RBLT<1> B_XWL<1> B_RWL<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<16> A_BLC_BOT<1> A_RBLC<1> A_BLT_BOT<1> A_RBLT<1> A_XWL<0> A_RWL<0> 
+ B_BLC_BOT<1> B_RBLC<1> B_BLT_BOT<1> B_RBLT<1> B_XWL<0> B_RWL<0> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<15> A_BLC_TOP<0> A_LBLC<15> A_BLT_TOP<0> A_LBLT<15> A_LWL<15> A_XWL<15> 
+ B_BLC_TOP<0> B_LBLC<15> B_BLT_TOP<0> B_LBLT<15> B_LWL<15> B_XWL<15> 
+ VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<14> A_LBLC<14> A_LBLC<15> A_LBLT<14> A_LBLT<15> A_LWL<14> A_XWL<14> 
+ B_LBLC<14> B_LBLC<15> B_LBLT<14> B_LBLT<15> B_LWL<14> B_XWL<14> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<13> A_LBLC<14> A_LBLC<13> A_LBLT<14> A_LBLT<13> A_LWL<13> A_XWL<13> 
+ B_LBLC<14> B_LBLC<13> B_LBLT<14> B_LBLT<13> B_LWL<13> B_XWL<13> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<12> A_LBLC<12> A_LBLC<13> A_LBLT<12> A_LBLT<13> A_LWL<12> A_XWL<12> 
+ B_LBLC<12> B_LBLC<13> B_LBLT<12> B_LBLT<13> B_LWL<12> B_XWL<12> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<11> A_LBLC<12> A_LBLC<11> A_LBLT<12> A_LBLT<11> A_LWL<11> A_XWL<11> 
+ B_LBLC<12> B_LBLC<11> B_LBLT<12> B_LBLT<11> B_LWL<11> B_XWL<11> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<10> A_LBLC<10> A_LBLC<11> A_LBLT<10> A_LBLT<11> A_LWL<10> A_XWL<10> 
+ B_LBLC<10> B_LBLC<11> B_LBLT<10> B_LBLT<11> B_LWL<10> B_XWL<10> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<9> A_LBLC<10> A_LBLC<9> A_LBLT<10> A_LBLT<9> A_LWL<9> A_XWL<9> 
+ B_LBLC<10> B_LBLC<9> B_LBLT<10> B_LBLT<9> B_LWL<9> B_XWL<9> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<8> A_LBLC<8> A_LBLC<9> A_LBLT<8> A_LBLT<9> A_LWL<8> A_XWL<8> B_LBLC<8> 
+ B_LBLC<9> B_LBLT<8> B_LBLT<9> B_LWL<8> B_XWL<8> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<7> A_LBLC<8> A_LBLC<7> A_LBLT<8> A_LBLT<7> A_LWL<7> A_XWL<7> B_LBLC<8> 
+ B_LBLC<7> B_LBLT<8> B_LBLT<7> B_LWL<7> B_XWL<7> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<6> A_LBLC<6> A_LBLC<7> A_LBLT<6> A_LBLT<7> A_LWL<6> A_XWL<6> B_LBLC<6> 
+ B_LBLC<7> B_LBLT<6> B_LBLT<7> B_LWL<6> B_XWL<6> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<5> A_LBLC<6> A_LBLC<5> A_LBLT<6> A_LBLT<5> A_LWL<5> A_XWL<5> B_LBLC<6> 
+ B_LBLC<5> B_LBLT<6> B_LBLT<5> B_LWL<5> B_XWL<5> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<4> A_LBLC<4> A_LBLC<5> A_LBLT<4> A_LBLT<5> A_LWL<4> A_XWL<4> B_LBLC<4> 
+ B_LBLC<5> B_LBLT<4> B_LBLT<5> B_LWL<4> B_XWL<4> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<3> A_LBLC<4> A_LBLC<3> A_LBLT<4> A_LBLT<3> A_LWL<3> A_XWL<3> B_LBLC<4> 
+ B_LBLC<3> B_LBLT<4> B_LBLT<3> B_LWL<3> B_XWL<3> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<2> A_LBLC<2> A_LBLC<3> A_LBLT<2> A_LBLT<3> A_LWL<2> A_XWL<2> B_LBLC<2> 
+ B_LBLC<3> B_LBLT<2> B_LBLT<3> B_LWL<2> B_XWL<2> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<1> A_LBLC<2> A_LBLC<1> A_LBLT<2> A_LBLT<1> A_LWL<1> A_XWL<1> B_LBLC<2> 
+ B_LBLC<1> B_LBLT<2> B_LBLT<1> B_LWL<1> B_XWL<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
XCELL<0> A_BLC_BOT<0> A_LBLC<1> A_BLT_BOT<0> A_LBLT<1> A_LWL<0> A_XWL<0> 
+ B_BLC_BOT<0> B_LBLC<1> B_BLT_BOT<0> B_LBLT<1> B_LWL<0> B_XWL<0> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_CELL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB A_BLC A_BLT B_BLC B_BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_16x2_EDGE_TB A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ B_BLC<1> B_BLC<0> B_BLT<1> B_BLT<0> VDD_CORE VSS
XEDGE<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB
XEDGE<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_TAP A_BLC A_BLT B_BLC B_BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_16x2_TAP A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ B_BLC<1> B_BLC<0> B_BLT<1> B_BLT<0> VDD_CORE VSS
XIEDGEBP_COL1<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL1<0> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL2<1> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL2<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_EDGE_TB
XITAP<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_TAP
XITAP<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_1024x64_c2_2P_BITKIT_TAP
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_TAP_LR NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BITKIT_16x2_TAP_LR VDD_CORE VSS
XCORNER<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER
XCORNER<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER
XTAP_BORDER VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_TAP_LR
.ENDS

.SUBCKT RSC_IHPSG13_CBUFX12 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=4.23u l=130.00n ng=6 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=9.72u l=130.00n ng=6 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDRV13X12 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX12 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=9.72u l=130.00n ng=6 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_WLDRV16X12 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX12
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_DEC04 ADDR<3> ADDR<2> ADDR<1> ADDR<0> CS ECLK_H_BOT 
+ ECLK_H_TOP ECLK_L_BOT ECLK_L_TOP WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> 
+ WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> VDD VSS
XI0<3> PADR<1> PADR<0> sel01<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<2> PADR<1> NADR<0> sel01<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<1> NADR<1> PADR<0> sel01<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<0> NADR<1> NADR<0> sel01<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI4 ECLK_L_BOT EN VDD VSS / RSC_IHPSG13_CINVX4
XI5 ECLK_H_BOT ECLK_L_BOT VDD VSS / RSC_IHPSG13_CINVX2
XI3<3> PADR<3> NADR<3> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> PADR<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> PADR<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> PADR<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XR0 ECLK_H_BOT ECLK_H_TOP / RSC_IHPSG13_MET2RES
XI11 ECLK_L_BOT ECLK_L_TOP / RSC_IHPSG13_MET2RES
XI1<3> PADR<2> PADR<3> CS sel23<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<2> PADR<3> CS sel23<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<2> NADR<3> CS sel23<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<2> NADR<3> CS sel23<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI2<15> sel23<3> sel01<3> EN WL<15> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<14> sel23<3> sel01<2> EN WL<14> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<13> sel23<3> sel01<1> EN WL<13> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<12> sel23<3> sel01<0> EN WL<12> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<11> sel23<2> sel01<3> EN WL<11> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<10> sel23<2> sel01<2> EN WL<10> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<9> sel23<2> sel01<1> EN WL<9> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<8> sel23<2> sel01<0> EN WL<8> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<7> sel23<1> sel01<3> EN WL<7> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<6> sel23<1> sel01<2> EN WL<6> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<5> sel23<1> sel01<1> EN WL<5> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<4> sel23<1> sel01<0> EN WL<4> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<3> sel23<0> sel01<3> EN WL<3> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<2> sel23<0> sel01<2> EN WL<2> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<1> sel23<0> sel01<1> EN WL<1> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<0> sel23<0> sel01<0> EN WL<0> VDD VSS / RSC_IHPSG13_NOR3X2
XCAPS4 VDD VSS / RSC_IHPSG13_FILLCAP4
XLATCH<3> CS ADDR<3> PADR<3> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<2> CS ADDR<2> PADR<2> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<1> CS ADDR<1> PADR<1> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<0> CS ADDR<0> PADR<0> VDD VSS / RSC_IHPSG13_LHPQX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_DEC02 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC ADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI2<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI2<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_DEC01 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC NADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI2<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI2<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_DEC00 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC NADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV<1> ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XADDRINV<0> ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_DEC03 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC ADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWDEC9 ADDR_N_I<8> ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> 
+ ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I 
+ WL_O<511> WL_O<510> WL_O<509> WL_O<508> WL_O<507> WL_O<506> WL_O<505> 
+ WL_O<504> WL_O<503> WL_O<502> WL_O<501> WL_O<500> WL_O<499> WL_O<498> 
+ WL_O<497> WL_O<496> WL_O<495> WL_O<494> WL_O<493> WL_O<492> WL_O<491> 
+ WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> WL_O<484> 
+ WL_O<483> WL_O<482> WL_O<481> WL_O<480> WL_O<479> WL_O<478> WL_O<477> 
+ WL_O<476> WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> 
+ WL_O<469> WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> WL_O<463> 
+ WL_O<462> WL_O<461> WL_O<460> WL_O<459> WL_O<458> WL_O<457> WL_O<456> 
+ WL_O<455> WL_O<454> WL_O<453> WL_O<452> WL_O<451> WL_O<450> WL_O<449> 
+ WL_O<448> WL_O<447> WL_O<446> WL_O<445> WL_O<444> WL_O<443> WL_O<442> 
+ WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> WL_O<436> WL_O<435> 
+ WL_O<434> WL_O<433> WL_O<432> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> WL_O<415> WL_O<414> 
+ WL_O<413> WL_O<412> WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> 
+ WL_O<406> WL_O<405> WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> 
+ WL_O<399> WL_O<398> WL_O<397> WL_O<396> WL_O<395> WL_O<394> WL_O<393> 
+ WL_O<392> WL_O<391> WL_O<390> WL_O<389> WL_O<388> WL_O<387> WL_O<386> 
+ WL_O<385> WL_O<384> WL_O<383> WL_O<382> WL_O<381> WL_O<380> WL_O<379> 
+ WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> WL_O<372> 
+ WL_O<371> WL_O<370> WL_O<369> WL_O<368> WL_O<367> WL_O<366> WL_O<365> 
+ WL_O<364> WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> 
+ WL_O<357> WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> WL_O<351> 
+ WL_O<350> WL_O<349> WL_O<348> WL_O<347> WL_O<346> WL_O<345> WL_O<344> 
+ WL_O<343> WL_O<342> WL_O<341> WL_O<340> WL_O<339> WL_O<338> WL_O<337> 
+ WL_O<336> WL_O<335> WL_O<334> WL_O<333> WL_O<332> WL_O<331> WL_O<330> 
+ WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> WL_O<324> WL_O<323> 
+ WL_O<322> WL_O<321> WL_O<320> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> WL_O<303> WL_O<302> 
+ WL_O<301> WL_O<300> WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> 
+ WL_O<294> WL_O<293> WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> 
+ WL_O<287> WL_O<286> WL_O<285> WL_O<284> WL_O<283> WL_O<282> WL_O<281> 
+ WL_O<280> WL_O<279> WL_O<278> WL_O<277> WL_O<276> WL_O<275> WL_O<274> 
+ WL_O<273> WL_O<272> WL_O<271> WL_O<270> WL_O<269> WL_O<268> WL_O<267> 
+ WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> WL_O<260> 
+ WL_O<259> WL_O<258> WL_O<257> WL_O<256> WL_O<255> WL_O<254> WL_O<253> 
+ WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> 
+ WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> WL_O<239> 
+ WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> WL_O<233> WL_O<232> 
+ WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> WL_O<226> WL_O<225> 
+ WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> WL_O<219> WL_O<218> 
+ WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> WL_O<212> WL_O<211> 
+ WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> WL_O<191> WL_O<190> 
+ WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> 
+ WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> 
+ WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> WL_O<170> WL_O<169> 
+ WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> WL_O<163> WL_O<162> 
+ WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> WL_O<156> WL_O<155> 
+ WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> WL_O<148> 
+ WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> WL_O<142> WL_O<141> 
+ WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> 
+ WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> WL_O<127> 
+ WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> 
+ WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> 
+ WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> 
+ WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> 
+ WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XSEL<31> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<31> ECLK_H<31> 
+ ECLK_H<32> ECLK_B<31> ECLK_B<32> WL_O<511> WL_O<510> WL_O<509> WL_O<508> 
+ WL_O<507> WL_O<506> WL_O<505> WL_O<504> WL_O<503> WL_O<502> WL_O<501> 
+ WL_O<500> WL_O<499> WL_O<498> WL_O<497> WL_O<496> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<30> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<30> ECLK_H<30> 
+ ECLK_H<31> ECLK_B<30> ECLK_B<31> WL_O<495> WL_O<494> WL_O<493> WL_O<492> 
+ WL_O<491> WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> 
+ WL_O<484> WL_O<483> WL_O<482> WL_O<481> WL_O<480> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<29> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<29> ECLK_H<29> 
+ ECLK_H<30> ECLK_B<29> ECLK_B<30> WL_O<479> WL_O<478> WL_O<477> WL_O<476> 
+ WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> WL_O<469> 
+ WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<28> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<28> ECLK_H<28> 
+ ECLK_H<29> ECLK_B<28> ECLK_B<29> WL_O<463> WL_O<462> WL_O<461> WL_O<460> 
+ WL_O<459> WL_O<458> WL_O<457> WL_O<456> WL_O<455> WL_O<454> WL_O<453> 
+ WL_O<452> WL_O<451> WL_O<450> WL_O<449> WL_O<448> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<27> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<27> ECLK_H<27> 
+ ECLK_H<28> ECLK_B<27> ECLK_B<28> WL_O<447> WL_O<446> WL_O<445> WL_O<444> 
+ WL_O<443> WL_O<442> WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> 
+ WL_O<436> WL_O<435> WL_O<434> WL_O<433> WL_O<432> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<26> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<26> ECLK_H<26> 
+ ECLK_H<27> ECLK_B<26> ECLK_B<27> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<25> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<25> ECLK_H<25> 
+ ECLK_H<26> ECLK_B<25> ECLK_B<26> WL_O<415> WL_O<414> WL_O<413> WL_O<412> 
+ WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> WL_O<406> WL_O<405> 
+ WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<24> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<24> ECLK_H<24> 
+ ECLK_H<25> ECLK_B<24> ECLK_B<25> WL_O<399> WL_O<398> WL_O<397> WL_O<396> 
+ WL_O<395> WL_O<394> WL_O<393> WL_O<392> WL_O<391> WL_O<390> WL_O<389> 
+ WL_O<388> WL_O<387> WL_O<386> WL_O<385> WL_O<384> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<23> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<23> ECLK_H<23> 
+ ECLK_H<24> ECLK_B<23> ECLK_B<24> WL_O<383> WL_O<382> WL_O<381> WL_O<380> 
+ WL_O<379> WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> 
+ WL_O<372> WL_O<371> WL_O<370> WL_O<369> WL_O<368> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<22> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<22> ECLK_H<22> 
+ ECLK_H<23> ECLK_B<22> ECLK_B<23> WL_O<367> WL_O<366> WL_O<365> WL_O<364> 
+ WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> WL_O<357> 
+ WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<21> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<21> ECLK_H<21> 
+ ECLK_H<22> ECLK_B<21> ECLK_B<22> WL_O<351> WL_O<350> WL_O<349> WL_O<348> 
+ WL_O<347> WL_O<346> WL_O<345> WL_O<344> WL_O<343> WL_O<342> WL_O<341> 
+ WL_O<340> WL_O<339> WL_O<338> WL_O<337> WL_O<336> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<20> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<20> ECLK_H<20> 
+ ECLK_H<21> ECLK_B<20> ECLK_B<21> WL_O<335> WL_O<334> WL_O<333> WL_O<332> 
+ WL_O<331> WL_O<330> WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> 
+ WL_O<324> WL_O<323> WL_O<322> WL_O<321> WL_O<320> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<19> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<19> ECLK_H<19> 
+ ECLK_H<20> ECLK_B<19> ECLK_B<20> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<18> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<18> ECLK_H<18> 
+ ECLK_H<19> ECLK_B<18> ECLK_B<19> WL_O<303> WL_O<302> WL_O<301> WL_O<300> 
+ WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> WL_O<294> WL_O<293> 
+ WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<17> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<17> ECLK_H<17> 
+ ECLK_H<18> ECLK_B<17> ECLK_B<18> WL_O<287> WL_O<286> WL_O<285> WL_O<284> 
+ WL_O<283> WL_O<282> WL_O<281> WL_O<280> WL_O<279> WL_O<278> WL_O<277> 
+ WL_O<276> WL_O<275> WL_O<274> WL_O<273> WL_O<272> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<16> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<16> ECLK_H<16> 
+ ECLK_H<17> ECLK_B<16> ECLK_B<17> WL_O<271> WL_O<270> WL_O<269> WL_O<268> 
+ WL_O<267> WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> 
+ WL_O<260> WL_O<259> WL_O<258> WL_O<257> WL_O<256> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XDEC10<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<30> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<26> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<22> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<18> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC01<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<29> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<25> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<21> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<17> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XL2<258> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<257> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<256> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<255> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<254> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<253> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<252> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<251> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<250> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<249> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<248> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<247> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<246> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<245> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<244> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<243> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<242> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<241> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<240> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<239> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<238> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<237> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<236> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<235> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<234> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<233> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<232> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<231> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<230> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<229> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<228> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<227> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<226> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<225> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<224> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<223> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<222> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<221> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<220> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<219> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<218> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<217> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<216> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<215> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<214> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<213> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<212> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<211> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<210> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<209> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<208> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<207> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<206> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<205> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<204> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<203> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<202> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<201> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<200> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<199> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<198> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<197> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<196> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<195> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<194> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<193> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<192> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<191> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<190> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<189> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<188> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<187> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<186> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<185> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<184> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<183> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<182> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<181> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<180> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<179> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<178> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<177> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<176> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<175> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<174> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<173> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<172> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<171> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<170> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<169> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<168> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<167> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<166> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<165> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<164> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<163> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<162> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<161> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<160> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<159> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<158> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<157> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<156> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<155> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<154> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<153> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<152> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<151> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<150> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<149> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<148> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<147> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<146> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<145> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<144> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<143> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<142> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<141> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<140> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<139> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<138> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<137> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<136> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<135> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<134> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<133> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC00<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<28> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<24> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<20> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<16> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC11<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<31> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<27> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<23> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<19> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XI0 ADDR_N_I<9> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWREG9 ACLK_N_I ADDR_I<8> ADDR_I<7> ADDR_I<6> ADDR_I<5> 
+ ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<8> ADDR_N_O<7> 
+ ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> 
+ ADDR_N_O<0> BIST_ADDR_I<8> BIST_ADDR_I<7> BIST_ADDR_I<6> BIST_ADDR_I<5> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XDFF<8> BIST_EN_I BIST_ADDR_I<8> ACLK_N_I ADDR_I<8> q_int<8> net04<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net04<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net04<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net04<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net04<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net04<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net04<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net04<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net04<8> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDRV<8> qn_int<8> ADDR_N_O<8> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XINV<8> q_int<8> qn_int<8> VDD VSS / RSC_IHPSG13_CINVX2
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_2P_DLY_MUX A SEL Z VDD VSS
XI11 net4 Z VDD VSS / RSC_IHPSG13_CINVX2
XI8 A D<3> SEL net4 VDD VSS / RSC_IHPSG13_MX2IX1
XI20<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_CTRL ACLK_N BIST_CK_I BIST_CS_I BIST_EN BIST_RE_I 
+ BIST_WE_I B_TIEL_O CK_I CS_I DCLK ECLK PULSE_H PULSE_L PULSE_O RCLK RE_I 
+ ROW_CS WCLK WE_I VDD VSS
XI17 ck_regs we col_we VDD VSS / RSC_IHPSG13_DFNQX2
XI16 ck_regs re col_re VDD VSS / RSC_IHPSG13_DFNQX2
XI18 ck_regs cs net7 VDD VSS / RSC_IHPSG13_DFNQX2
XI71 ACLK_N net012 PULSE_O VDD VSS / RSC_IHPSG13_DFNQX2
XI77 col_we net017 net016 VDD VSS / RSC_IHPSG13_CNAND2X2
XI76 col_re net017 net018 VDD VSS / RSC_IHPSG13_CNAND2X2
XI15 ck_dly WEorREandCS aclk VDD VSS / RSC_IHPSG13_CGATEPX4
XI14 ck WEandCS DCLK VDD VSS / RSC_IHPSG13_CGATEPX4
XI60 net7 ROW_CS VDD VSS / RSC_IHPSG13_CBUFX8
XI73 PULSE_O net012 VDD VSS / RSC_IHPSG13_CINVX2
XI8 net017 net8 VDD VSS / RSC_IHPSG13_CINVX2
XCAPS4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XBM_TIEL B_TIEL_O VDD VSS / RSC_IHPSG13_TIEL
XI64 ck ck_dly VDD VSS / RSC_IHPSG13_CDLYX2
XI86 CS_I BIST_CS_I BIST_EN cs VDD VSS / RSC_IHPSG13_MX2X2
XI87 CK_I BIST_CK_I BIST_EN ck VDD VSS / RSC_IHPSG13_MX2X2
XI85 WE_I BIST_WE_I BIST_EN we VDD VSS / RSC_IHPSG13_MX2X2
XI84 RE_I BIST_RE_I BIST_EN re VDD VSS / RSC_IHPSG13_MX2X2
XI48 ck_dly ck_regs VDD VSS / RSC_IHPSG13_CINVX4
XI81 net016 WCLK VDD VSS / RSC_IHPSG13_CINVX4
XI80 net018 RCLK VDD VSS / RSC_IHPSG13_CINVX4
XI78 net8 net020 VDD VSS / RSC_IHPSG13_CINVX4
XCAPS8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI6 PULSE_L PULSE_H net017 VDD VSS / RSC_IHPSG13_XOR2X2
XI22 we cs WEandCS VDD VSS / RSC_IHPSG13_AND2X2
XI79 net020 ECLK VDD VSS / RSC_IHPSG13_CINVX8
XI63 aclk ACLK_N VDD VSS / RSC_IHPSG13_CINVX8
XI21 re we cs WEorREandCS VDD VSS / RSC_IHPSG13_OA12X1
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDEC5 ACLK_N ADDR<4> ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<4> BIST_ADDR<3> 
+ BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<4> BIST_EN_I BIST_ADDR<4> ACLK_N ADDR<4> addr_int<1> net13<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int<0> net13<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net13<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net13<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net13<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI15<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI15<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> addr_int<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_CBUFX2
XI13<0> addr_int<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XI14<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_BLDRV A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> 
+ A_SEL_P<1> A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> 
+ B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> 
+ B_SEL_P<2> B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS
MA_CWN<3> A_BLC<3> A_BLC_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<2> A_BLC<2> A_BLC_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<1> A_BLC<1> A_BLC_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<0> A_BLC<0> A_BLC_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<3> A_BLT<3> A_BLT_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<2> A_BLT<2> A_BLT_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<1> A_BLT<1> A_BLT_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<0> A_BLT<0> A_BLT_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<3> B_BLT<3> B_BLT_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<2> B_BLT<2> B_BLT_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<1> B_BLT<1> B_BLT_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<0> B_BLT<0> B_BLT_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<3> B_BLC<3> B_BLC_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<2> B_BLC<2> B_BLC_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<1> B_BLC<1> B_BLC_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<0> B_BLC<0> B_BLC_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CPR<3> A_BLC<3> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<2> A_BLC<2> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<1> A_BLC<1> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<0> A_BLC<0> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TWP<3> A_BLT<3> A_BLT_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<2> A_BLT<2> A_BLT_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<1> A_BLT<1> A_BLT_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<0> A_BLT<0> A_BLT_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<3> A_BLC<3> A_BLC_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<2> A_BLC<2> A_BLC_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<1> A_BLC<1> A_BLC_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<0> A_BLC<0> A_BLC_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TPR<3> A_BLT<3> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<2> A_BLT<2> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<1> A_BLT<1> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<0> A_BLT<0> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TSP<3> A_BLT_SEL A_SEL_N<3> A_BLT<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<2> A_BLT_SEL A_SEL_N<2> A_BLT<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<1> A_BLT_SEL A_SEL_N<1> A_BLT<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<0> A_BLT_SEL A_SEL_N<0> A_BLT<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<3> A_BLC_SEL A_SEL_N<3> A_BLC<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<2> A_BLC_SEL A_SEL_N<2> A_BLC<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<1> A_BLC_SEL A_SEL_N<1> A_BLC<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<0> A_BLC_SEL A_SEL_N<0> A_BLC<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<3> B_BLC<3> B_BLC_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<2> B_BLC<2> B_BLC_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<1> B_BLC<1> B_BLC_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<0> B_BLC<0> B_BLC_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<3> B_BLT<3> B_BLT_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<2> B_BLT<2> B_BLT_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<1> B_BLT<1> B_BLT_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<0> B_BLT<0> B_BLT_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<3> B_BLT_SEL B_SEL_N<3> B_BLT<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<2> B_BLT_SEL B_SEL_N<2> B_BLT<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<1> B_BLT_SEL B_SEL_N<1> B_BLT<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<0> B_BLT_SEL B_SEL_N<0> B_BLT<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TPR<3> B_BLT<3> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<2> B_BLT<2> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<1> B_BLT<1> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<0> B_BLT<0> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CSP<3> B_BLC_SEL B_SEL_N<3> B_BLC<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<2> B_BLC_SEL B_SEL_N<2> B_BLC<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<1> B_BLC_SEL B_SEL_N<1> B_BLC<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<0> B_BLC_SEL B_SEL_N<0> B_BLC<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CPR<3> B_BLC<3> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<2> B_BLC<2> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<1> B_BLC<1> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<0> B_BLC<0> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
XA_SEL<3> A_SEL_P<3> A_SEL_N<3> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<2> A_SEL_P<2> A_SEL_N<2> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<1> A_SEL_P<1> A_SEL_N<1> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<0> A_SEL_P<0> A_SEL_N<0> VDD VSS / RSC_IHPSG13_INVX2
XA_CINV<3> A_BLT_PMOS_DRIVE<3> A_BLC_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<2> A_BLT_PMOS_DRIVE<2> A_BLC_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<1> A_BLT_PMOS_DRIVE<1> A_BLC_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<0> A_BLT_PMOS_DRIVE<0> A_BLC_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<3> A_BLC_PMOS_DRIVE<3> A_BLT_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<2> A_BLC_PMOS_DRIVE<2> A_BLT_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<1> A_BLC_PMOS_DRIVE<1> A_BLT_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<0> A_BLC_PMOS_DRIVE<0> A_BLT_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_SEL<3> B_SEL_P<3> B_SEL_N<3> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<2> B_SEL_P<2> B_SEL_N<2> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<1> B_SEL_P<1> B_SEL_N<1> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<0> B_SEL_P<0> B_SEL_N<0> VDD VSS / RSC_IHPSG13_INVX2
XB_TINV<3> B_BLC_PMOS_DRIVE<3> B_BLT_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<2> B_BLC_PMOS_DRIVE<2> B_BLT_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<1> B_BLC_PMOS_DRIVE<1> B_BLT_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<0> B_BLC_PMOS_DRIVE<0> B_BLT_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<3> B_BLT_PMOS_DRIVE<3> B_BLC_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<2> B_BLT_PMOS_DRIVE<2> B_BLC_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<1> B_BLT_PMOS_DRIVE<1> B_BLC_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<0> B_BLT_PMOS_DRIVE<0> B_BLC_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TDEC<3> A_SEL_P<3> A_WR_ONE A_BLT_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<2> A_SEL_P<2> A_WR_ONE A_BLT_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<1> A_SEL_P<1> A_WR_ONE A_BLT_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<0> A_SEL_P<0> A_WR_ONE A_BLT_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<3> A_SEL_P<3> A_WR_ZERO A_BLC_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<2> A_SEL_P<2> A_WR_ZERO A_BLC_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<1> A_SEL_P<1> A_WR_ZERO A_BLC_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<0> A_SEL_P<0> A_WR_ZERO A_BLC_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<3> B_SEL_P<3> B_WR_ZERO B_BLC_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<2> B_SEL_P<2> B_WR_ZERO B_BLC_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<1> B_SEL_P<1> B_WR_ZERO B_BLC_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<0> B_SEL_P<0> B_WR_ZERO B_BLC_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<3> B_SEL_P<3> B_WR_ONE B_BLT_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<2> B_SEL_P<2> B_WR_ONE B_BLT_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<1> B_SEL_P<1> B_WR_ONE B_BLT_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<0> B_SEL_P<0> B_WR_ONE B_BLT_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
.ENDS
.SUBCKT RSC_IHPSG13_AND2X6 A B Z VDD VSS
MN3 Z net6 VSS VSS nmos m=1 w=2.94u l=130.00n ng=3 nrd=0 nrs=0
MN4 net9 B VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD pmos m=1 w=4.86u l=130.00n ng=3 nrd=0 nrs=0
MP0 net6 B VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLCTRL5 A_ADDR_COL<1> A_ADDR_COL<0> A_ADDR_DEC<7> 
+ A_ADDR_DEC<6> A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<31> 
+ A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> 
+ A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> 
+ A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> 
+ A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> 
+ A_BLC<1> A_BLC<0> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> 
+ A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> 
+ A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> 
+ A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_COL<1> B_ADDR_COL<0> 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> 
+ B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I 
+ B_BIST_EN_I B_BLC<31> B_BLC<30> B_BLC<29> B_BLC<28> B_BLC<27> B_BLC<26> 
+ B_BLC<25> B_BLC<24> B_BLC<23> B_BLC<22> B_BLC<21> B_BLC<20> B_BLC<19> 
+ B_BLC<18> B_BLC<17> B_BLC<16> B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> 
+ B_BLC<11> B_BLC<10> B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> 
+ B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<31> B_BLT<30> B_BLT<29> B_BLT<28> 
+ B_BLT<27> B_BLT<26> B_BLT<25> B_BLT<24> B_BLT<23> B_BLT<22> B_BLT<21> 
+ B_BLT<20> B_BLT<19> B_BLT<18> B_BLT<17> B_BLT<16> B_BLT<15> B_BLT<14> 
+ B_BLT<13> B_BLT<12> B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> 
+ B_BLT<5> B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L 
+ B_DCLK_B_R B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L 
+ B_RCLK_R B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_I80<1> B_WCLK_B_L B_RCLK_B_L B_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XB_I80<0> B_WCLK_B_L B_RCLK_B_L B_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<1> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<0> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XI_FILL4<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XB_INV<6> B_N1<1> B_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<5> B_N0<1> B_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<4> B_N0<0> B_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<3> B_ADDR_COL<1> B_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<2> B_ADDR_COL<1> B_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<1> B_ADDR_COL<0> B_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<0> B_ADDR_COL<0> B_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<6> A_N1<1> A_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<5> A_N0<1> A_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<4> A_N0<0> A_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<3> A_ADDR_COL<1> A_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<2> A_ADDR_COL<1> A_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_ADDR_COL<0> A_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL<0> A_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_I81<3> B_W_nor_R<1> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<2> B_W_nor_R<1> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<1> B_W_nor_R<0> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<0> B_W_nor_R<0> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<3> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<2> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XI_FILL8<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XAB_BLMUX<7> A_BLC<31> A_BLC<30> A_BLC<29> A_BLC<28> A_BLC_SEL A_BLT<31> 
+ A_BLT<30> A_BLT<29> A_BLT<28> A_BLT_SEL A_PRE_N A_SEL_P<31> A_SEL_P<30> 
+ A_SEL_P<29> A_SEL_P<28> A_WR_ONE A_WR_ZERO B_BLC<31> B_BLC<30> B_BLC<29> 
+ B_BLC<28> B_BLC_SEL B_BLT<31> B_BLT<30> B_BLT<29> B_BLT<28> B_BLT_SEL 
+ B_PRE_N B_SEL_P<31> B_SEL_P<30> B_SEL_P<29> B_SEL_P<28> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<6> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> A_BLC_SEL A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT_SEL A_PRE_N A_SEL_P<27> A_SEL_P<26> 
+ A_SEL_P<25> A_SEL_P<24> A_WR_ONE A_WR_ZERO B_BLC<27> B_BLC<26> B_BLC<25> 
+ B_BLC<24> B_BLC_SEL B_BLT<27> B_BLT<26> B_BLT<25> B_BLT<24> B_BLT_SEL 
+ B_PRE_N B_SEL_P<27> B_SEL_P<26> B_SEL_P<25> B_SEL_P<24> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<5> A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC_SEL A_BLT<23> 
+ A_BLT<22> A_BLT<21> A_BLT<20> A_BLT_SEL A_PRE_N A_SEL_P<23> A_SEL_P<22> 
+ A_SEL_P<21> A_SEL_P<20> A_WR_ONE A_WR_ZERO B_BLC<23> B_BLC<22> B_BLC<21> 
+ B_BLC<20> B_BLC_SEL B_BLT<23> B_BLT<22> B_BLT<21> B_BLT<20> B_BLT_SEL 
+ B_PRE_N B_SEL_P<23> B_SEL_P<22> B_SEL_P<21> B_SEL_P<20> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<4> A_BLC<19> A_BLC<18> A_BLC<17> A_BLC<16> A_BLC_SEL A_BLT<19> 
+ A_BLT<18> A_BLT<17> A_BLT<16> A_BLT_SEL A_PRE_N A_SEL_P<19> A_SEL_P<18> 
+ A_SEL_P<17> A_SEL_P<16> A_WR_ONE A_WR_ZERO B_BLC<19> B_BLC<18> B_BLC<17> 
+ B_BLC<16> B_BLC_SEL B_BLT<19> B_BLT<18> B_BLT<17> B_BLT<16> B_BLT_SEL 
+ B_PRE_N B_SEL_P<19> B_SEL_P<18> B_SEL_P<17> B_SEL_P<16> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<3> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC_SEL A_BLT<15> 
+ A_BLT<14> A_BLT<13> A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<15> A_SEL_P<14> 
+ A_SEL_P<13> A_SEL_P<12> A_WR_ONE A_WR_ZERO B_BLC<15> B_BLC<14> B_BLC<13> 
+ B_BLC<12> B_BLC_SEL B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT_SEL 
+ B_PRE_N B_SEL_P<15> B_SEL_P<14> B_SEL_P<13> B_SEL_P<12> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<2> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC_SEL A_BLT<11> 
+ A_BLT<10> A_BLT<9> A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<11> A_SEL_P<10> 
+ A_SEL_P<9> A_SEL_P<8> A_WR_ONE A_WR_ZERO B_BLC<11> B_BLC<10> B_BLC<9> 
+ B_BLC<8> B_BLC_SEL B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT_SEL B_PRE_N 
+ B_SEL_P<11> B_SEL_P<10> B_SEL_P<9> B_SEL_P<8> B_WR_ONE B_WR_ZERO VDD 
+ VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<7> A_SEL_P<6> A_SEL_P<5> 
+ A_SEL_P<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC_SEL 
+ B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N B_SEL_P<7> B_SEL_P<6> 
+ B_SEL_P<5> B_SEL_P<4> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> A_SEL_P<1> 
+ A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLC_SEL 
+ B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> B_SEL_P<2> 
+ B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BLDRV
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<31> net041<0> B_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<30> net041<1> B_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<29> net041<2> B_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<28> net041<3> B_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<27> net041<4> B_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<26> net041<5> B_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<25> net041<6> B_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<24> net041<7> B_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<23> net041<8> B_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<22> net041<9> B_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<21> net041<10> B_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<20> net041<11> B_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<19> net041<12> B_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<18> net041<13> B_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<17> net041<14> B_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<16> net041<15> B_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<15> net041<16> B_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<14> net041<17> B_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<13> net041<18> B_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<12> net041<19> B_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<11> net041<20> B_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<10> net041<21> B_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<9> net041<22> B_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<8> net041<23> B_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<7> net041<24> B_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<6> net041<25> B_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<5> net041<26> B_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<4> net041<27> B_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<3> net041<28> B_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<2> net041<29> B_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<1> net041<30> B_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<0> net041<31> B_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<31> net23<0> A_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<30> net23<1> A_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<29> net23<2> A_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<28> net23<3> A_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<27> net23<4> A_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<26> net23<5> A_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<25> net23<6> A_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<24> net23<7> A_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<23> net23<8> A_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<22> net23<9> A_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<21> net23<10> A_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<20> net23<11> A_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<19> net23<12> A_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<18> net23<13> A_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<17> net23<14> A_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<16> net23<15> A_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<15> net23<16> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<17> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<18> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<19> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<20> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<21> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<22> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<23> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<24> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<25> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<26> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<27> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<28> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<29> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<30> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<31> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net042 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net043 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net21 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_DEC3<31> B_P1<1> B_P0<1> B_ADDR_DEC<7> net041<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<30> B_P1<1> B_P0<1> B_ADDR_DEC<6> net041<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<29> B_P1<1> B_P0<1> B_ADDR_DEC<5> net041<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<28> B_P1<1> B_P0<1> B_ADDR_DEC<4> net041<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<27> B_P1<1> B_P0<1> B_ADDR_DEC<3> net041<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<26> B_P1<1> B_P0<1> B_ADDR_DEC<2> net041<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<25> B_P1<1> B_P0<1> B_ADDR_DEC<1> net041<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<24> B_P1<1> B_P0<1> B_ADDR_DEC<0> net041<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<23> B_P1<1> B_N0<1> B_ADDR_DEC<7> net041<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<22> B_P1<1> B_N0<1> B_ADDR_DEC<6> net041<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<21> B_P1<1> B_N0<1> B_ADDR_DEC<5> net041<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<20> B_P1<1> B_N0<1> B_ADDR_DEC<4> net041<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<19> B_P1<1> B_N0<1> B_ADDR_DEC<3> net041<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<18> B_P1<1> B_N0<1> B_ADDR_DEC<2> net041<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<17> B_P1<1> B_N0<1> B_ADDR_DEC<1> net041<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<16> B_P1<1> B_N0<1> B_ADDR_DEC<0> net041<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<15> B_N1<0> B_P0<0> B_ADDR_DEC<7> net041<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<14> B_N1<0> B_P0<0> B_ADDR_DEC<6> net041<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<13> B_N1<0> B_P0<0> B_ADDR_DEC<5> net041<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<12> B_N1<0> B_P0<0> B_ADDR_DEC<4> net041<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<11> B_N1<0> B_P0<0> B_ADDR_DEC<3> net041<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<10> B_N1<0> B_P0<0> B_ADDR_DEC<2> net041<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<9> B_N1<0> B_P0<0> B_ADDR_DEC<1> net041<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<8> B_N1<0> B_P0<0> B_ADDR_DEC<0> net041<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<7> B_N1<0> B_N0<0> B_ADDR_DEC<7> net041<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<6> B_N1<0> B_N0<0> B_ADDR_DEC<6> net041<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<5> B_N1<0> B_N0<0> B_ADDR_DEC<5> net041<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<4> B_N1<0> B_N0<0> B_ADDR_DEC<4> net041<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<3> B_N1<0> B_N0<0> B_ADDR_DEC<3> net041<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<2> B_N1<0> B_N0<0> B_ADDR_DEC<2> net041<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<1> B_N1<0> B_N0<0> B_ADDR_DEC<1> net041<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<0> B_N1<0> B_N0<0> B_ADDR_DEC<0> net041<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<31> A_P1<1> A_P0<1> A_ADDR_DEC<7> net23<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<30> A_P1<1> A_P0<1> A_ADDR_DEC<6> net23<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<29> A_P1<1> A_P0<1> A_ADDR_DEC<5> net23<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<28> A_P1<1> A_P0<1> A_ADDR_DEC<4> net23<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<27> A_P1<1> A_P0<1> A_ADDR_DEC<3> net23<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<26> A_P1<1> A_P0<1> A_ADDR_DEC<2> net23<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<25> A_P1<1> A_P0<1> A_ADDR_DEC<1> net23<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<24> A_P1<1> A_P0<1> A_ADDR_DEC<0> net23<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<23> A_P1<1> A_N0<1> A_ADDR_DEC<7> net23<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<22> A_P1<1> A_N0<1> A_ADDR_DEC<6> net23<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<21> A_P1<1> A_N0<1> A_ADDR_DEC<5> net23<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<20> A_P1<1> A_N0<1> A_ADDR_DEC<4> net23<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<19> A_P1<1> A_N0<1> A_ADDR_DEC<3> net23<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<18> A_P1<1> A_N0<1> A_ADDR_DEC<2> net23<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<17> A_P1<1> A_N0<1> A_ADDR_DEC<1> net23<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<16> A_P1<1> A_N0<1> A_ADDR_DEC<0> net23<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<15> A_N1<0> A_P0<0> A_ADDR_DEC<7> net23<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<14> A_N1<0> A_P0<0> A_ADDR_DEC<6> net23<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<13> A_N1<0> A_P0<0> A_ADDR_DEC<5> net23<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<12> A_N1<0> A_P0<0> A_ADDR_DEC<4> net23<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<11> A_N1<0> A_P0<0> A_ADDR_DEC<3> net23<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<10> A_N1<0> A_P0<0> A_ADDR_DEC<2> net23<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<9> A_N1<0> A_P0<0> A_ADDR_DEC<1> net23<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<8> A_N1<0> A_P0<0> A_ADDR_DEC<0> net23<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<7> A_N1<0> A_N0<0> A_ADDR_DEC<7> net23<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<6> A_N1<0> A_N0<0> A_ADDR_DEC<6> net23<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<5> A_N1<0> A_N0<0> A_ADDR_DEC<5> net23<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<4> A_N1<0> A_N0<0> A_ADDR_DEC<4> net23<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<3> A_N1<0> A_N0<0> A_ADDR_DEC<3> net23<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<2> A_N1<0> A_N0<0> A_ADDR_DEC<2> net23<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<1> A_N1<0> A_N0<0> A_ADDR_DEC<1> net23<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<0> A_N1<0> A_N0<0> A_ADDR_DEC<0> net23<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDRV13_FILL4 VDD VSS
XI0<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RSC_IHPSG13_CBUFX16 A Z VDD VSS
MN0 net4 A VSS VSS nmos m=1 w=2.115u l=130.00n ng=3 nrd=0 nrs=0
MN1 Z net4 VSS VSS nmos m=1 w=5.64u l=130.00n ng=8 nrd=0 nrs=0
MP1 Z net4 VDD VDD pmos m=1 w=13.000u l=130.00n ng=8 nrd=0 
+ nrs=0
MP0 net4 A VDD VDD pmos m=1 w=4.89u l=130.00n ng=3 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDRV13X16 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX16 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=12.96u l=130.00n ng=8 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_WLDRV16X16 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX16
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDRV13X4 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1 VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_WLDRV16X4 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWDEC8 ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> 
+ ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<255> 
+ WL_O<254> WL_O<253> WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> 
+ WL_O<247> WL_O<246> WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> 
+ WL_O<240> WL_O<239> WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> 
+ WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> 
+ WL_O<226> WL_O<225> WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> 
+ WL_O<205> WL_O<204> WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> 
+ WL_O<198> WL_O<197> WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> 
+ WL_O<191> WL_O<190> WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> 
+ WL_O<184> WL_O<183> WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> 
+ WL_O<177> WL_O<176> WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> 
+ WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> 
+ WL_O<163> WL_O<162> WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> 
+ WL_O<156> WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> 
+ WL_O<149> WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> 
+ WL_O<142> WL_O<141> WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> 
+ WL_O<135> WL_O<134> WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> 
+ WL_O<128> WL_O<127> WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> 
+ WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> 
+ WL_O<114> WL_O<113> WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> 
+ WL_O<92> WL_O<91> WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> 
+ WL_O<84> WL_O<83> WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> 
+ WL_O<76> WL_O<75> WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> 
+ WL_O<68> WL_O<67> WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> 
+ WL_O<60> WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> 
+ WL_O<52> WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> 
+ WL_O<44> WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> 
+ WL_O<36> WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> 
+ WL_O<28> WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> 
+ WL_O<20> WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> 
+ WL_O<12> WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> 
+ WL_O<3> WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XDEC10<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC00<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC01<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWREG8 ACLK_N_I ADDR_I<7> ADDR_I<6> ADDR_I<5> ADDR_I<4> 
+ ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<7> ADDR_N_O<6> ADDR_N_O<5> 
+ ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<7> 
+ BIST_ADDR_I<6> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> 
+ BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI10 VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDEC4 ACLK_N ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<3> BIST_ADDR<2> 
+ BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int net12<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net12<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net12<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net12<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI14 addr_int ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI15 ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLCTRL4 A_ADDR_COL A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<15> A_BLC<14> 
+ A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> 
+ A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> 
+ A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L 
+ A_DCLK_B_R A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L 
+ A_RCLK_R A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_COL 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> 
+ B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I 
+ B_BIST_EN_I B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> B_BLC<11> B_BLC<10> 
+ B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC<3> B_BLC<2> 
+ B_BLC<1> B_BLC<0> B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT<11> 
+ B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT<3> 
+ B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L B_DCLK_B_R B_DCLK_L B_DCLK_R 
+ B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L B_RCLK_R B_TIEH_O B_WCLK_B_L 
+ B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_I80 B_RCLK_B_L B_WCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_RCLK_B_L A_WCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XI_FILL4<26> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<25> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<24> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<23> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<22> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<21> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<20> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<19> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<18> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<17> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<1> B_N0 B_P0 VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<0> B_ADDR_COL B_N0 VDD VSS / RSC_IHPSG13_CINVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_N0 A_P0 VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL A_N0 VDD VSS / RSC_IHPSG13_CINVX4
XB_I81<1> net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<0> net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XAB_BLMUX<3> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC_SEL A_BLT<15> 
+ A_BLT<14> A_BLT<13> A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<15> A_SEL_P<14> 
+ A_SEL_P<13> A_SEL_P<12> A_WR_ONE A_WR_ZERO B_BLC<15> B_BLC<14> B_BLC<13> 
+ B_BLC<12> B_BLC_SEL B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT_SEL 
+ B_PRE_N B_SEL_P<15> B_SEL_P<14> B_SEL_P<13> B_SEL_P<12> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<2> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC_SEL A_BLT<11> 
+ A_BLT<10> A_BLT<9> A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<11> A_SEL_P<10> 
+ A_SEL_P<9> A_SEL_P<8> A_WR_ONE A_WR_ZERO B_BLC<11> B_BLC<10> B_BLC<9> 
+ B_BLC<8> B_BLC_SEL B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT_SEL B_PRE_N 
+ B_SEL_P<11> B_SEL_P<10> B_SEL_P<9> B_SEL_P<8> B_WR_ONE B_WR_ZERO VDD 
+ VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<7> A_SEL_P<6> A_SEL_P<5> 
+ A_SEL_P<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC_SEL 
+ B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N B_SEL_P<7> B_SEL_P<6> 
+ B_SEL_P<5> B_SEL_P<4> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> A_SEL_P<1> 
+ A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLC_SEL 
+ B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> B_SEL_P<2> 
+ B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_BLDRV
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net046 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net045 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net24 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3INV<15> net23<0> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<1> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<2> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<3> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<4> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<5> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<6> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<7> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<8> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<9> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<10> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<11> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<12> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<13> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<14> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<15> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<15> net044<0> B_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<14> net044<1> B_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<13> net044<2> B_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<12> net044<3> B_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<11> net044<4> B_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<10> net044<5> B_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<9> net044<6> B_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<8> net044<7> B_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<7> net044<8> B_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<6> net044<9> B_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<5> net044<10> B_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<4> net044<11> B_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<3> net044<12> B_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<2> net044<13> B_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<1> net044<14> B_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<0> net044<15> B_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XI_FILL8<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_DEC3<15> A_P0 A_ADDR_DEC<7> net23<0> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<14> A_P0 A_ADDR_DEC<6> net23<1> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<13> A_P0 A_ADDR_DEC<5> net23<2> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<12> A_P0 A_ADDR_DEC<4> net23<3> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<11> A_P0 A_ADDR_DEC<3> net23<4> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<10> A_P0 A_ADDR_DEC<2> net23<5> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<9> A_P0 A_ADDR_DEC<1> net23<6> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<8> A_P0 A_ADDR_DEC<0> net23<7> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<7> A_N0 A_ADDR_DEC<7> net23<8> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<6> A_N0 A_ADDR_DEC<6> net23<9> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<5> A_N0 A_ADDR_DEC<5> net23<10> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<4> A_N0 A_ADDR_DEC<4> net23<11> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<3> A_N0 A_ADDR_DEC<3> net23<12> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<2> A_N0 A_ADDR_DEC<2> net23<13> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<1> A_N0 A_ADDR_DEC<1> net23<14> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<0> A_N0 A_ADDR_DEC<0> net23<15> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<15> B_P0 B_ADDR_DEC<7> net044<0> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<14> B_P0 B_ADDR_DEC<6> net044<1> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<13> B_P0 B_ADDR_DEC<5> net044<2> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<12> B_P0 B_ADDR_DEC<4> net044<3> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<11> B_P0 B_ADDR_DEC<3> net044<4> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<10> B_P0 B_ADDR_DEC<2> net044<5> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<9> B_P0 B_ADDR_DEC<1> net044<6> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<8> B_P0 B_ADDR_DEC<0> net044<7> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<7> B_N0 B_ADDR_DEC<7> net044<8> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<6> B_N0 B_ADDR_DEC<6> net044<9> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<5> B_N0 B_ADDR_DEC<5> net044<10> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<4> B_N0 B_ADDR_DEC<4> net044<11> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<3> B_N0 B_ADDR_DEC<3> net044<12> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<2> B_N0 B_ADDR_DEC<2> net044<13> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<1> B_N0 B_ADDR_DEC<1> net044<14> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<0> B_N0 B_ADDR_DEC<0> net044<15> VDD VSS / RSC_IHPSG13_NAND2X2
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWDEC5 ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> 
+ ADDR_N_I<0> CS_I ECLK_I WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0 ADDR_N_I<5> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWREG5 ACLK_N_I ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> 
+ ADDR_I<0> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDEC3 ACLK_N ADDR<2> ADDR<1> ADDR<0> ADDR_COL<1> 
+ ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> 
+ ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> 
+ BIST_EN_I VDD VSS
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net13<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net13<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net13<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_DFPQD_MSAFFX2P CP DN DP QN QP VDD VSS
XI_AMP CP DN DP QN QP VDD VSS / RSC_IHPSG13_DFPQD_MSAFFX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLCTRL3 A_ADDR_DEC<7> A_ADDR_DEC<6> A_ADDR_DEC<5> 
+ A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> A_ADDR_DEC<0> 
+ A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> 
+ A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R A_DCLK_L 
+ A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R A_TIEH_O 
+ A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_DEC<7> B_ADDR_DEC<6> 
+ B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> 
+ B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I B_BIST_EN_I B_BLC<7> B_BLC<6> B_BLC<5> 
+ B_BLC<4> B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<7> B_BLT<6> B_BLT<5> 
+ B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L B_DCLK_B_R 
+ B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L B_RCLK_R 
+ B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net044 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net043 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2P
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2P
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> 
+ B_BLC<4> B_BLC_SEL B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> 
+ B_BLC<0> B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I80 B_WCLK_B_L B_RCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DO_WRITE_P B_DI_N B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XB_I75 B_DO_WRITE_P B_DI_R B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_WCLK_B_L A_RCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XB_I81 net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWDEC6 ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> 
+ ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<63> WL_O<62> WL_O<61> WL_O<60> 
+ WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> 
+ WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> 
+ WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> 
+ WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> 
+ WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> 
+ WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> 
+ WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> 
+ WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC10 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XDEC11 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWREG6 ACLK_N_I ADDR_I<5> ADDR_I<4> ADDR_I<3> ADDR_I<2> 
+ ADDR_I<1> ADDR_I<0> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> 
+ ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDRV13X16 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XI1<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_WLDRV16X16 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX16
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_DEC01 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC NADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XI2 VDD VSS / RSC_IHPSG13_FILLCAP4
XADDRINV ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_DEC00 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC NADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV<1> ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XADDRINV<0> ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1 VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWDEC5 ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> 
+ ADDR_N_I<0> CS_I ECLK_I WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XI0 ADDR_N_I<5> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWREG5 ACLK_N_I ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> 
+ ADDR_I<0> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDEC5 ACLK_N ADDR<4> ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<4> BIST_ADDR<3> 
+ BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<1> addr_int<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_CBUFX2
XI13<0> addr_int<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XDFF<4> BIST_EN_I BIST_ADDR<4> ACLK_N ADDR<4> addr_int<1> net7<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int<0> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net7<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI15<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI15<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLCTRL5 A_ADDR_COL<1> A_ADDR_COL<0> A_ADDR_DEC<7> 
+ A_ADDR_DEC<6> A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<31> 
+ A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> 
+ A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> 
+ A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> 
+ A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> 
+ A_BLC<1> A_BLC<0> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> 
+ A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> 
+ A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> 
+ A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_I80<1> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<0> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XI80<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_INV<6> A_N1<1> A_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<5> A_N0<1> A_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<4> A_N0<0> A_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<3> A_ADDR_COL<1> A_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<2> A_ADDR_COL<1> A_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_ADDR_COL<0> A_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL<0> A_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_I81<3> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<2> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<31> A_BLC<31> A_BLC_SEL A_BLT<31> A_BLT_SEL A_PRE_N A_SEL_P<31> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<30> A_BLC<30> A_BLC_SEL A_BLT<30> A_BLT_SEL A_PRE_N A_SEL_P<30> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<29> A_BLC<29> A_BLC_SEL A_BLT<29> A_BLT_SEL A_PRE_N A_SEL_P<29> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<28> A_BLC<28> A_BLC_SEL A_BLT<28> A_BLT_SEL A_PRE_N A_SEL_P<28> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<27> A_BLC<27> A_BLC_SEL A_BLT<27> A_BLT_SEL A_PRE_N A_SEL_P<27> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<26> A_BLC<26> A_BLC_SEL A_BLT<26> A_BLT_SEL A_PRE_N A_SEL_P<26> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<25> A_BLC<25> A_BLC_SEL A_BLT<25> A_BLT_SEL A_PRE_N A_SEL_P<25> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<24> A_BLC<24> A_BLC_SEL A_BLT<24> A_BLT_SEL A_PRE_N A_SEL_P<24> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<23> A_BLC<23> A_BLC_SEL A_BLT<23> A_BLT_SEL A_PRE_N A_SEL_P<23> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<22> A_BLC<22> A_BLC_SEL A_BLT<22> A_BLT_SEL A_PRE_N A_SEL_P<22> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<21> A_BLC<21> A_BLC_SEL A_BLT<21> A_BLT_SEL A_PRE_N A_SEL_P<21> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<20> A_BLC<20> A_BLC_SEL A_BLT<20> A_BLT_SEL A_PRE_N A_SEL_P<20> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<19> A_BLC<19> A_BLC_SEL A_BLT<19> A_BLT_SEL A_PRE_N A_SEL_P<19> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<18> A_BLC<18> A_BLC_SEL A_BLT<18> A_BLT_SEL A_PRE_N A_SEL_P<18> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<17> A_BLC<17> A_BLC_SEL A_BLT<17> A_BLT_SEL A_PRE_N A_SEL_P<17> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<16> A_BLC<16> A_BLC_SEL A_BLT<16> A_BLT_SEL A_PRE_N A_SEL_P<16> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<15> A_BLC<15> A_BLC_SEL A_BLT<15> A_BLT_SEL A_PRE_N A_SEL_P<15> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<14> A_BLC<14> A_BLC_SEL A_BLT<14> A_BLT_SEL A_PRE_N A_SEL_P<14> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<13> A_BLC<13> A_BLC_SEL A_BLT<13> A_BLT_SEL A_PRE_N A_SEL_P<13> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<12> A_BLC<12> A_BLC_SEL A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<12> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<11> A_BLC<11> A_BLC_SEL A_BLT<11> A_BLT_SEL A_PRE_N A_SEL_P<11> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<10> A_BLC<10> A_BLC_SEL A_BLT<10> A_BLT_SEL A_PRE_N A_SEL_P<10> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<9> A_BLC<9> A_BLC_SEL A_BLT<9> A_BLT_SEL A_PRE_N A_SEL_P<9> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<8> A_BLC<8> A_BLC_SEL A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<8> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_SEL_P<7> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_SEL_P<6> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_SEL_P<5> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<4> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_SEL_P<3> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_SEL_P<2> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_SEL_P<1> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<0> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_1024x64_c2_1P_BLDRV
XA_CAPS<17> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<31> net23<0> A_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<30> net23<1> A_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<29> net23<2> A_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<28> net23<3> A_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<27> net23<4> A_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<26> net23<5> A_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<25> net23<6> A_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<24> net23<7> A_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<23> net23<8> A_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<22> net23<9> A_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<21> net23<10> A_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<20> net23<11> A_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<19> net23<12> A_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<18> net23<13> A_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<17> net23<14> A_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<16> net23<15> A_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<15> net23<16> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<17> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<18> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<19> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<20> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<21> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<22> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<23> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<24> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<25> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<26> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<27> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<28> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<29> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<30> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<31> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net21 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3<31> A_P1<1> A_P0<1> A_ADDR_DEC<7> net23<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<30> A_P1<1> A_P0<1> A_ADDR_DEC<6> net23<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<29> A_P1<1> A_P0<1> A_ADDR_DEC<5> net23<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<28> A_P1<1> A_P0<1> A_ADDR_DEC<4> net23<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<27> A_P1<1> A_P0<1> A_ADDR_DEC<3> net23<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<26> A_P1<1> A_P0<1> A_ADDR_DEC<2> net23<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<25> A_P1<1> A_P0<1> A_ADDR_DEC<1> net23<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<24> A_P1<1> A_P0<1> A_ADDR_DEC<0> net23<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<23> A_P1<1> A_N0<1> A_ADDR_DEC<7> net23<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<22> A_P1<1> A_N0<1> A_ADDR_DEC<6> net23<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<21> A_P1<1> A_N0<1> A_ADDR_DEC<5> net23<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<20> A_P1<1> A_N0<1> A_ADDR_DEC<4> net23<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<19> A_P1<1> A_N0<1> A_ADDR_DEC<3> net23<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<18> A_P1<1> A_N0<1> A_ADDR_DEC<2> net23<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<17> A_P1<1> A_N0<1> A_ADDR_DEC<1> net23<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<16> A_P1<1> A_N0<1> A_ADDR_DEC<0> net23<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<15> A_N1<0> A_P0<0> A_ADDR_DEC<7> net23<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<14> A_N1<0> A_P0<0> A_ADDR_DEC<6> net23<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<13> A_N1<0> A_P0<0> A_ADDR_DEC<5> net23<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<12> A_N1<0> A_P0<0> A_ADDR_DEC<4> net23<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<11> A_N1<0> A_P0<0> A_ADDR_DEC<3> net23<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<10> A_N1<0> A_P0<0> A_ADDR_DEC<2> net23<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<9> A_N1<0> A_P0<0> A_ADDR_DEC<1> net23<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<8> A_N1<0> A_P0<0> A_ADDR_DEC<0> net23<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<7> A_N1<0> A_N0<0> A_ADDR_DEC<7> net23<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<6> A_N1<0> A_N0<0> A_ADDR_DEC<6> net23<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<5> A_N1<0> A_N0<0> A_ADDR_DEC<5> net23<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<4> A_N1<0> A_N0<0> A_ADDR_DEC<4> net23<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<3> A_N1<0> A_N0<0> A_ADDR_DEC<3> net23<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<2> A_N1<0> A_N0<0> A_ADDR_DEC<2> net23<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<1> A_N1<0> A_N0<0> A_ADDR_DEC<1> net23<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<0> A_N1<0> A_N0<0> A_ADDR_DEC<0> net23<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDRV13X12 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_WLDRV16X12 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX12
.ENDS



.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDRV13X8 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX8 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_WLDRV16X8 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX8
.ENDS



.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDEC2 ACLK_N ADDR<1> ADDR<0> ADDR_COL<1> ADDR_COL<0> 
+ ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> ADDR_DEC<2> 
+ ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI16<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<3> PADR<0> PADR<1> addr_n<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<2> NADR<0> PADR<1> addr_n<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<1> PADR<0> NADR<1> addr_n<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<0> NADR<0> NADR<1> addr_n<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI17<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI17<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI14<3> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_TIEL
XI14<2> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_TIEL
XI14<1> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_TIEL
XI14<0> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_TIEL
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net12<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net12<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI15<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLCTRL2 A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<3> A_BLC<2> A_BLC<1> 
+ A_BLC<0> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_DEC<3> B_ADDR_DEC<2> 
+ B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I B_BIST_EN_I B_BLC<3> 
+ B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I 
+ B_DCLK_B_L B_DCLK_B_R B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R 
+ B_RCLK_L B_RCLK_R B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD 
+ VSS
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net046 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net045 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_CAPS VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS VDD VSS / RSC_IHPSG13_FILLCAP4
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XB_I80 B_RCLK_B_L B_WCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_RCLK_B_L A_WCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XB_I44 B_WCLK_B_L B_BM_N B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_WCLK_B_L A_BM_N A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_I81 net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XAB_BLMUX A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> 
+ B_BLC<0> B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_1024x64_c2_2P_BLDRV
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net039 net040 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_I51 net039 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_COLDRV13_FILL4C2 VDD VSS
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWDEC7 ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> 
+ ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<127> WL_O<126> 
+ WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> 
+ WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> 
+ WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> WL_O<105> 
+ WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> WL_O<98> WL_O<97> 
+ WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> WL_O<90> WL_O<89> 
+ WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> WL_O<82> WL_O<81> 
+ WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> WL_O<74> WL_O<73> 
+ WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> WL_O<66> WL_O<65> 
+ WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> WL_O<58> WL_O<57> 
+ WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> WL_O<50> WL_O<49> 
+ WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> WL_O<42> WL_O<41> 
+ WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> WL_O<34> WL_O<33> 
+ WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> WL_O<26> WL_O<25> 
+ WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> WL_O<18> WL_O<17> 
+ WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC03
XDEC01<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC01
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC02
XDEC00<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_2P_DEC00
XI0 ADDR_N_I<7> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWREG7 ACLK_N_I ADDR_I<6> ADDR_I<5> ADDR_I<4> ADDR_I<3> 
+ ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<6> 
+ BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> 
+ BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWDEC4 ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> 
+ CS_I ECLK_I WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XSEL ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I ECLK_H<1> 
+ ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> 
+ WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> 
+ WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_2P_DEC04
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_2P_ROWREG4 ACLK_N_I ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net7<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_TAP BLC BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_TAP A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ VDD_CORE VSS
XITAP<1> A_BLC<1> A_BLT<1> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_1P_BITKIT_TAP
XITAP<0> A_BLC<0> A_BLT<0> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_1024x64_c2_1P_BITKIT_TAP
XIEDGEBP_COL1<1> BLC<1> BLT<1> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL1<0> BLC<1> BLT<1> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL2<1> BLC<0> BLT<0> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL2<0> BLC<0> BLT<0> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_EDGE_TB
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_TAP_LR VDD_CORE VSS
XCORNER<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER
XCORNER<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_CORNER
XTAP_BORDER VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_1024x64_c2_1P_BITKIT_TAP_LR
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_DEC03 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI0 VDD VSS / RSC_IHPSG13_FILLCAP4
XDEC ADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_DEC02 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC ADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XI2 VDD VSS / RSC_IHPSG13_FILLCAP4
XADDRINV ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWDEC8 ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> 
+ ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<255> 
+ WL_O<254> WL_O<253> WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> 
+ WL_O<247> WL_O<246> WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> 
+ WL_O<240> WL_O<239> WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> 
+ WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> 
+ WL_O<226> WL_O<225> WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> 
+ WL_O<205> WL_O<204> WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> 
+ WL_O<198> WL_O<197> WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> 
+ WL_O<191> WL_O<190> WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> 
+ WL_O<184> WL_O<183> WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> 
+ WL_O<177> WL_O<176> WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> 
+ WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> 
+ WL_O<163> WL_O<162> WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> 
+ WL_O<156> WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> 
+ WL_O<149> WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> 
+ WL_O<142> WL_O<141> WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> 
+ WL_O<135> WL_O<134> WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> 
+ WL_O<128> WL_O<127> WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> 
+ WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> 
+ WL_O<114> WL_O<113> WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> 
+ WL_O<92> WL_O<91> WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> 
+ WL_O<84> WL_O<83> WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> 
+ WL_O<76> WL_O<75> WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> 
+ WL_O<68> WL_O<67> WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> 
+ WL_O<60> WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> 
+ WL_O<52> WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> 
+ WL_O<44> WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> 
+ WL_O<36> WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> 
+ WL_O<28> WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> 
+ WL_O<20> WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> 
+ WL_O<12> WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> 
+ WL_O<3> WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC10<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC00<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XDEC01<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWREG8 ACLK_N_I ADDR_I<7> ADDR_I<6> ADDR_I<5> ADDR_I<4> 
+ ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<7> ADDR_N_O<6> ADDR_N_O<5> 
+ ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<7> 
+ BIST_ADDR_I<6> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> 
+ BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWDEC9 ADDR_N_I<8> ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> 
+ ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I 
+ WL_O<511> WL_O<510> WL_O<509> WL_O<508> WL_O<507> WL_O<506> WL_O<505> 
+ WL_O<504> WL_O<503> WL_O<502> WL_O<501> WL_O<500> WL_O<499> WL_O<498> 
+ WL_O<497> WL_O<496> WL_O<495> WL_O<494> WL_O<493> WL_O<492> WL_O<491> 
+ WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> WL_O<484> 
+ WL_O<483> WL_O<482> WL_O<481> WL_O<480> WL_O<479> WL_O<478> WL_O<477> 
+ WL_O<476> WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> 
+ WL_O<469> WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> WL_O<463> 
+ WL_O<462> WL_O<461> WL_O<460> WL_O<459> WL_O<458> WL_O<457> WL_O<456> 
+ WL_O<455> WL_O<454> WL_O<453> WL_O<452> WL_O<451> WL_O<450> WL_O<449> 
+ WL_O<448> WL_O<447> WL_O<446> WL_O<445> WL_O<444> WL_O<443> WL_O<442> 
+ WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> WL_O<436> WL_O<435> 
+ WL_O<434> WL_O<433> WL_O<432> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> WL_O<415> WL_O<414> 
+ WL_O<413> WL_O<412> WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> 
+ WL_O<406> WL_O<405> WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> 
+ WL_O<399> WL_O<398> WL_O<397> WL_O<396> WL_O<395> WL_O<394> WL_O<393> 
+ WL_O<392> WL_O<391> WL_O<390> WL_O<389> WL_O<388> WL_O<387> WL_O<386> 
+ WL_O<385> WL_O<384> WL_O<383> WL_O<382> WL_O<381> WL_O<380> WL_O<379> 
+ WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> WL_O<372> 
+ WL_O<371> WL_O<370> WL_O<369> WL_O<368> WL_O<367> WL_O<366> WL_O<365> 
+ WL_O<364> WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> 
+ WL_O<357> WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> WL_O<351> 
+ WL_O<350> WL_O<349> WL_O<348> WL_O<347> WL_O<346> WL_O<345> WL_O<344> 
+ WL_O<343> WL_O<342> WL_O<341> WL_O<340> WL_O<339> WL_O<338> WL_O<337> 
+ WL_O<336> WL_O<335> WL_O<334> WL_O<333> WL_O<332> WL_O<331> WL_O<330> 
+ WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> WL_O<324> WL_O<323> 
+ WL_O<322> WL_O<321> WL_O<320> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> WL_O<303> WL_O<302> 
+ WL_O<301> WL_O<300> WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> 
+ WL_O<294> WL_O<293> WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> 
+ WL_O<287> WL_O<286> WL_O<285> WL_O<284> WL_O<283> WL_O<282> WL_O<281> 
+ WL_O<280> WL_O<279> WL_O<278> WL_O<277> WL_O<276> WL_O<275> WL_O<274> 
+ WL_O<273> WL_O<272> WL_O<271> WL_O<270> WL_O<269> WL_O<268> WL_O<267> 
+ WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> WL_O<260> 
+ WL_O<259> WL_O<258> WL_O<257> WL_O<256> WL_O<255> WL_O<254> WL_O<253> 
+ WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> 
+ WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> WL_O<239> 
+ WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> WL_O<233> WL_O<232> 
+ WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> WL_O<226> WL_O<225> 
+ WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> WL_O<219> WL_O<218> 
+ WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> WL_O<212> WL_O<211> 
+ WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> WL_O<191> WL_O<190> 
+ WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> 
+ WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> 
+ WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> WL_O<170> WL_O<169> 
+ WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> WL_O<163> WL_O<162> 
+ WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> WL_O<156> WL_O<155> 
+ WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> WL_O<148> 
+ WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> WL_O<142> WL_O<141> 
+ WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> 
+ WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> WL_O<127> 
+ WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> 
+ WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> 
+ WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> 
+ WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> 
+ WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XL2<172> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<171> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<170> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<169> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<168> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<167> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<166> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<165> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<164> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<163> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<162> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<161> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<160> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<159> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<158> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<157> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<156> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<155> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<154> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<153> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<152> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<151> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<150> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<149> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<148> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<147> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<146> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<145> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<144> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<143> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<142> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<141> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<140> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<139> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<138> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<137> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<136> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<135> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<134> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<133> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC11<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<31> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<27> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<23> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<19> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC00<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<28> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<24> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<20> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<16> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XSEL<31> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<31> ECLK_H<31> 
+ ECLK_H<32> ECLK_B<31> ECLK_B<32> WL_O<511> WL_O<510> WL_O<509> WL_O<508> 
+ WL_O<507> WL_O<506> WL_O<505> WL_O<504> WL_O<503> WL_O<502> WL_O<501> 
+ WL_O<500> WL_O<499> WL_O<498> WL_O<497> WL_O<496> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<30> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<30> ECLK_H<30> 
+ ECLK_H<31> ECLK_B<30> ECLK_B<31> WL_O<495> WL_O<494> WL_O<493> WL_O<492> 
+ WL_O<491> WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> 
+ WL_O<484> WL_O<483> WL_O<482> WL_O<481> WL_O<480> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<29> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<29> ECLK_H<29> 
+ ECLK_H<30> ECLK_B<29> ECLK_B<30> WL_O<479> WL_O<478> WL_O<477> WL_O<476> 
+ WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> WL_O<469> 
+ WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<28> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<28> ECLK_H<28> 
+ ECLK_H<29> ECLK_B<28> ECLK_B<29> WL_O<463> WL_O<462> WL_O<461> WL_O<460> 
+ WL_O<459> WL_O<458> WL_O<457> WL_O<456> WL_O<455> WL_O<454> WL_O<453> 
+ WL_O<452> WL_O<451> WL_O<450> WL_O<449> WL_O<448> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<27> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<27> ECLK_H<27> 
+ ECLK_H<28> ECLK_B<27> ECLK_B<28> WL_O<447> WL_O<446> WL_O<445> WL_O<444> 
+ WL_O<443> WL_O<442> WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> 
+ WL_O<436> WL_O<435> WL_O<434> WL_O<433> WL_O<432> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<26> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<26> ECLK_H<26> 
+ ECLK_H<27> ECLK_B<26> ECLK_B<27> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<25> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<25> ECLK_H<25> 
+ ECLK_H<26> ECLK_B<25> ECLK_B<26> WL_O<415> WL_O<414> WL_O<413> WL_O<412> 
+ WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> WL_O<406> WL_O<405> 
+ WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<24> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<24> ECLK_H<24> 
+ ECLK_H<25> ECLK_B<24> ECLK_B<25> WL_O<399> WL_O<398> WL_O<397> WL_O<396> 
+ WL_O<395> WL_O<394> WL_O<393> WL_O<392> WL_O<391> WL_O<390> WL_O<389> 
+ WL_O<388> WL_O<387> WL_O<386> WL_O<385> WL_O<384> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<23> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<23> ECLK_H<23> 
+ ECLK_H<24> ECLK_B<23> ECLK_B<24> WL_O<383> WL_O<382> WL_O<381> WL_O<380> 
+ WL_O<379> WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> 
+ WL_O<372> WL_O<371> WL_O<370> WL_O<369> WL_O<368> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<22> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<22> ECLK_H<22> 
+ ECLK_H<23> ECLK_B<22> ECLK_B<23> WL_O<367> WL_O<366> WL_O<365> WL_O<364> 
+ WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> WL_O<357> 
+ WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<21> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<21> ECLK_H<21> 
+ ECLK_H<22> ECLK_B<21> ECLK_B<22> WL_O<351> WL_O<350> WL_O<349> WL_O<348> 
+ WL_O<347> WL_O<346> WL_O<345> WL_O<344> WL_O<343> WL_O<342> WL_O<341> 
+ WL_O<340> WL_O<339> WL_O<338> WL_O<337> WL_O<336> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<20> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<20> ECLK_H<20> 
+ ECLK_H<21> ECLK_B<20> ECLK_B<21> WL_O<335> WL_O<334> WL_O<333> WL_O<332> 
+ WL_O<331> WL_O<330> WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> 
+ WL_O<324> WL_O<323> WL_O<322> WL_O<321> WL_O<320> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<19> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<19> ECLK_H<19> 
+ ECLK_H<20> ECLK_B<19> ECLK_B<20> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<18> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<18> ECLK_H<18> 
+ ECLK_H<19> ECLK_B<18> ECLK_B<19> WL_O<303> WL_O<302> WL_O<301> WL_O<300> 
+ WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> WL_O<294> WL_O<293> 
+ WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<17> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<17> ECLK_H<17> 
+ ECLK_H<18> ECLK_B<17> ECLK_B<18> WL_O<287> WL_O<286> WL_O<285> WL_O<284> 
+ WL_O<283> WL_O<282> WL_O<281> WL_O<280> WL_O<279> WL_O<278> WL_O<277> 
+ WL_O<276> WL_O<275> WL_O<274> WL_O<273> WL_O<272> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<16> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<16> ECLK_H<16> 
+ ECLK_H<17> ECLK_B<16> ECLK_B<17> WL_O<271> WL_O<270> WL_O<269> WL_O<268> 
+ WL_O<267> WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> 
+ WL_O<260> WL_O<259> WL_O<258> WL_O<257> WL_O<256> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XDEC01<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<29> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<25> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<21> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<17> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC10<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<30> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<26> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<22> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<18> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XI0 ADDR_N_I<9> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWREG9 ACLK_N_I ADDR_I<8> ADDR_I<7> ADDR_I<6> ADDR_I<5> 
+ ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<8> ADDR_N_O<7> 
+ ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> 
+ ADDR_N_O<0> BIST_ADDR_I<8> BIST_ADDR_I<7> BIST_ADDR_I<6> BIST_ADDR_I<5> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<8> q_int<8> qn_int<8> VDD VSS / RSC_IHPSG13_CINVX2
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<8> qn_int<8> ADDR_N_O<8> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<8> BIST_EN_I BIST_ADDR_I<8> ACLK_N_I ADDR_I<8> q_int<8> net04<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net04<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net04<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net04<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net04<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net04<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net04<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net04<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net04<8> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWDEC7 ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> 
+ ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<127> WL_O<126> 
+ WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> 
+ WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> 
+ WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> WL_O<105> 
+ WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> WL_O<98> WL_O<97> 
+ WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> WL_O<90> WL_O<89> 
+ WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> WL_O<82> WL_O<81> 
+ WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> WL_O<74> WL_O<73> 
+ WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> WL_O<66> WL_O<65> 
+ WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> WL_O<58> WL_O<57> 
+ WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> WL_O<50> WL_O<49> 
+ WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> WL_O<42> WL_O<41> 
+ WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> WL_O<34> WL_O<33> 
+ WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> WL_O<26> WL_O<25> 
+ WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> WL_O<18> WL_O<17> 
+ WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XDEC00<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC01<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0 ADDR_N_I<7> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWREG7 ACLK_N_I ADDR_I<6> ADDR_I<5> ADDR_I<4> ADDR_I<3> 
+ ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<6> 
+ BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> 
+ BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS

.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLDRV13X8 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_WLDRV16X8 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX8
.ENDS



.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWDEC6 ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> 
+ ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<63> WL_O<62> WL_O<61> WL_O<60> 
+ WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> 
+ WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> 
+ WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> 
+ WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> 
+ WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> 
+ WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> 
+ WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> 
+ WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<3> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC03
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC00
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC01
XDEC10 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<2> VDD VSS / 
+ RM_IHPSG13_1024x64_c2_1P_DEC02
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_1024x64_c2_1P_DEC04
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_1024x64_c2_1P_ROWREG6 ACLK_N_I ADDR_I<5> ADDR_I<4> ADDR_I<3> ADDR_I<2> 
+ ADDR_I<1> ADDR_I<0> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> 
+ ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0 A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<255> A_LWL<254> A_LWL<253> A_LWL<252> A_LWL<251> A_LWL<250> A_LWL<249> A_LWL<248> A_LWL<247> A_LWL<246> A_LWL<245> A_LWL<244> A_LWL<243> A_LWL<242> A_LWL<241> A_LWL<240> A_LWL<239> A_LWL<238> A_LWL<237> A_LWL<236> A_LWL<235> A_LWL<234> A_LWL<233> A_LWL<232> A_LWL<231> A_LWL<230> A_LWL<229> A_LWL<228> A_LWL<227> A_LWL<226> A_LWL<225> A_LWL<224> A_LWL<223> A_LWL<222> A_LWL<221> A_LWL<220> A_LWL<219> A_LWL<218> A_LWL<217> A_LWL<216> A_LWL<215> A_LWL<214> A_LWL<213> A_LWL<212> A_LWL<211> A_LWL<210> A_LWL<209> A_LWL<208> A_LWL<207> A_LWL<206> A_LWL<205> A_LWL<204> A_LWL<203> A_LWL<202> A_LWL<201> A_LWL<200> A_LWL<199> A_LWL<198> A_LWL<197> A_LWL<196> A_LWL<195> A_LWL<194> A_LWL<193> A_LWL<192> A_LWL<191> A_LWL<190> A_LWL<189> A_LWL<188> A_LWL<187> A_LWL<186> A_LWL<185> A_LWL<184> A_LWL<183> A_LWL<182> A_LWL<181> A_LWL<180> A_LWL<179> A_LWL<178> A_LWL<177> A_LWL<176> A_LWL<175> A_LWL<174> A_LWL<173> A_LWL<172> A_LWL<171> A_LWL<170> A_LWL<169> A_LWL<168> A_LWL<167> A_LWL<166> A_LWL<165> A_LWL<164> A_LWL<163> A_LWL<162> A_LWL<161> A_LWL<160> A_LWL<159> A_LWL<158> A_LWL<157> A_LWL<156> A_LWL<155> A_LWL<154> A_LWL<153> A_LWL<152> A_LWL<151> A_LWL<150> A_LWL<149> A_LWL<148> A_LWL<147> A_LWL<146> A_LWL<145> A_LWL<144> A_LWL<143> A_LWL<142> A_LWL<141> A_LWL<140> A_LWL<139> A_LWL<138> A_LWL<137> A_LWL<136> A_LWL<135> A_LWL<134> A_LWL<133> A_LWL<132> A_LWL<131> A_LWL<130> A_LWL<129> A_LWL<128> A_LWL<127> A_LWL<126> A_LWL<125> A_LWL<124> A_LWL<123> A_LWL<122> A_LWL<121> A_LWL<120> A_LWL<119> A_LWL<118> A_LWL<117> A_LWL<116> A_LWL<115> A_LWL<114> A_LWL<113> A_LWL<112> A_LWL<111> A_LWL<110> A_LWL<109> A_LWL<108> A_LWL<107> A_LWL<106> A_LWL<105> A_LWL<104> A_LWL<103> A_LWL<102> A_LWL<101> A_LWL<100> A_LWL<99> A_LWL<98> A_LWL<97> A_LWL<96> A_LWL<95> A_LWL<94> A_LWL<93> A_LWL<92> A_LWL<91> A_LWL<90> A_LWL<89> A_LWL<88> A_LWL<87> A_LWL<86> A_LWL<85> A_LWL<84> A_LWL<83> A_LWL<82> A_LWL<81> A_LWL<80> A_LWL<79> A_LWL<78> A_LWL<77> A_LWL<76> A_LWL<75> A_LWL<74> A_LWL<73> A_LWL<72> A_LWL<71> A_LWL<70> A_LWL<69> A_LWL<68> A_LWL<67> A_LWL<66> A_LWL<65> A_LWL<64> A_LWL<63> A_LWL<62> A_LWL<61> A_LWL<60> A_LWL<59> A_LWL<58> A_LWL<57> A_LWL<56> A_LWL<55> A_LWL<54> A_LWL<53> A_LWL<52> A_LWL<51> A_LWL<50> A_LWL<49> A_LWL<48> A_LWL<47> A_LWL<46> A_LWL<45> A_LWL<44> A_LWL<43> A_LWL<42> A_LWL<41> A_LWL<40> A_LWL<39> A_LWL<38> A_LWL<37> A_LWL<36> A_LWL<35> A_LWL<34> A_LWL<33> A_LWL<32> A_LWL<31> A_LWL<30> A_LWL<29> A_LWL<28> A_LWL<27> A_LWL<26> A_LWL<25> A_LWL<24> A_LWL<23> A_LWL<22> A_LWL<21> A_LWL<20> A_LWL<19> A_LWL<18> A_LWL<17> A_LWL<16> A_LWL<15> A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<255> A_RWL<254> A_RWL<253> A_RWL<252> A_RWL<251> A_RWL<250> A_RWL<249> A_RWL<248> A_RWL<247> A_RWL<246> A_RWL<245> A_RWL<244> A_RWL<243> A_RWL<242> A_RWL<241> A_RWL<240> A_RWL<239> A_RWL<238> A_RWL<237> A_RWL<236> A_RWL<235> A_RWL<234> A_RWL<233> A_RWL<232> A_RWL<231> A_RWL<230> A_RWL<229> A_RWL<228> A_RWL<227> A_RWL<226> A_RWL<225> A_RWL<224> A_RWL<223> A_RWL<222> A_RWL<221> A_RWL<220> A_RWL<219> A_RWL<218> A_RWL<217> A_RWL<216> A_RWL<215> A_RWL<214> A_RWL<213> A_RWL<212> A_RWL<211> A_RWL<210> A_RWL<209> A_RWL<208> A_RWL<207> A_RWL<206> A_RWL<205> A_RWL<204> A_RWL<203> A_RWL<202> A_RWL<201> A_RWL<200> A_RWL<199> A_RWL<198> A_RWL<197> A_RWL<196> A_RWL<195> A_RWL<194> A_RWL<193> A_RWL<192> A_RWL<191> A_RWL<190> A_RWL<189> A_RWL<188> A_RWL<187> A_RWL<186> A_RWL<185> A_RWL<184> A_RWL<183> A_RWL<182> A_RWL<181> A_RWL<180> A_RWL<179> A_RWL<178> A_RWL<177> A_RWL<176> A_RWL<175> A_RWL<174> A_RWL<173> A_RWL<172> A_RWL<171> A_RWL<170> A_RWL<169> A_RWL<168> A_RWL<167> A_RWL<166> A_RWL<165> A_RWL<164> A_RWL<163> A_RWL<162> A_RWL<161> A_RWL<160> A_RWL<159> A_RWL<158> A_RWL<157> A_RWL<156> A_RWL<155> A_RWL<154> A_RWL<153> A_RWL<152> A_RWL<151> A_RWL<150> A_RWL<149> A_RWL<148> A_RWL<147> A_RWL<146> A_RWL<145> A_RWL<144> A_RWL<143> A_RWL<142> A_RWL<141> A_RWL<140> A_RWL<139> A_RWL<138> A_RWL<137> A_RWL<136> A_RWL<135> A_RWL<134> A_RWL<133> A_RWL<132> A_RWL<131> A_RWL<130> A_RWL<129> A_RWL<128> A_RWL<127> A_RWL<126> A_RWL<125> A_RWL<124> A_RWL<123> A_RWL<122> A_RWL<121> A_RWL<120> A_RWL<119> A_RWL<118> A_RWL<117> A_RWL<116> A_RWL<115> A_RWL<114> A_RWL<113> A_RWL<112> A_RWL<111> A_RWL<110> A_RWL<109> A_RWL<108> A_RWL<107> A_RWL<106> A_RWL<105> A_RWL<104> A_RWL<103> A_RWL<102> A_RWL<101> A_RWL<100> A_RWL<99> A_RWL<98> A_RWL<97> A_RWL<96> A_RWL<95> A_RWL<94> A_RWL<93> A_RWL<92> A_RWL<91> A_RWL<90> A_RWL<89> A_RWL<88> A_RWL<87> A_RWL<86> A_RWL<85> A_RWL<84> A_RWL<83> A_RWL<82> A_RWL<81> A_RWL<80> A_RWL<79> A_RWL<78> A_RWL<77> A_RWL<76> A_RWL<75> A_RWL<74> A_RWL<73> A_RWL<72> A_RWL<71> A_RWL<70> A_RWL<69> A_RWL<68> A_RWL<67> A_RWL<66> A_RWL<65> A_RWL<64> A_RWL<63> A_RWL<62> A_RWL<61> A_RWL<60> A_RWL<59> A_RWL<58> A_RWL<57> A_RWL<56> A_RWL<55> A_RWL<54> A_RWL<53> A_RWL<52> A_RWL<51> A_RWL<50> A_RWL<49> A_RWL<48> A_RWL<47> A_RWL<46> A_RWL<45> A_RWL<44> A_RWL<43> A_RWL<42> A_RWL<41> A_RWL<40> A_RWL<39> A_RWL<38> A_RWL<37> A_RWL<36> A_RWL<35> A_RWL<34> A_RWL<33> A_RWL<32> A_RWL<31> A_RWL<30> A_RWL<29> A_RWL<28> A_RWL<27> A_RWL<26> A_RWL<25> A_RWL<24> A_RWL<23> A_RWL<22> A_RWL<21> A_RWL<20> A_RWL<19> A_RWL<18> A_RWL<17> A_RWL<16> A_RWL<15> A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE VSS
XRAM<16> A_BLC<29> A_BLC<28> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT<29> A_BLT<28> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<255> A_LWL<254> A_LWL<253> A_LWL<252> A_LWL<251> A_LWL<250> A_LWL<249> A_LWL<248> A_LWL<247> A_LWL<246> A_LWL<245> A_LWL<244> A_LWL<243> A_LWL<242> A_LWL<241> A_LWL<240> A_RWL<255> A_RWL<254> A_RWL<253> A_RWL<252> A_RWL<251> A_RWL<250> A_RWL<249> A_RWL<248> A_RWL<247> A_RWL<246> A_RWL<245> A_RWL<244> A_RWL<243> A_RWL<242> A_RWL<241> A_RWL<240> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<15> A_BLC<27> A_BLC<26> A_BLC<29> A_BLC<28> A_BLT<27> A_BLT<26> A_BLT<29> A_BLT<28> A_LWL<239> A_LWL<238> A_LWL<237> A_LWL<236> A_LWL<235> A_LWL<234> A_LWL<233> A_LWL<232> A_LWL<231> A_LWL<230> A_LWL<229> A_LWL<228> A_LWL<227> A_LWL<226> A_LWL<225> A_LWL<224> A_RWL<239> A_RWL<238> A_RWL<237> A_RWL<236> A_RWL<235> A_RWL<234> A_RWL<233> A_RWL<232> A_RWL<231> A_RWL<230> A_RWL<229> A_RWL<228> A_RWL<227> A_RWL<226> A_RWL<225> A_RWL<224> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<14> A_BLC<25> A_BLC<24> A_BLC<27> A_BLC<26> A_BLT<25> A_BLT<24> A_BLT<27> A_BLT<26> A_LWL<223> A_LWL<222> A_LWL<221> A_LWL<220> A_LWL<219> A_LWL<218> A_LWL<217> A_LWL<216> A_LWL<215> A_LWL<214> A_LWL<213> A_LWL<212> A_LWL<211> A_LWL<210> A_LWL<209> A_LWL<208> A_RWL<223> A_RWL<222> A_RWL<221> A_RWL<220> A_RWL<219> A_RWL<218> A_RWL<217> A_RWL<216> A_RWL<215> A_RWL<214> A_RWL<213> A_RWL<212> A_RWL<211> A_RWL<210> A_RWL<209> A_RWL<208> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<13> A_BLC<23> A_BLC<22> A_BLC<25> A_BLC<24> A_BLT<23> A_BLT<22> A_BLT<25> A_BLT<24> A_LWL<207> A_LWL<206> A_LWL<205> A_LWL<204> A_LWL<203> A_LWL<202> A_LWL<201> A_LWL<200> A_LWL<199> A_LWL<198> A_LWL<197> A_LWL<196> A_LWL<195> A_LWL<194> A_LWL<193> A_LWL<192> A_RWL<207> A_RWL<206> A_RWL<205> A_RWL<204> A_RWL<203> A_RWL<202> A_RWL<201> A_RWL<200> A_RWL<199> A_RWL<198> A_RWL<197> A_RWL<196> A_RWL<195> A_RWL<194> A_RWL<193> A_RWL<192> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<12> A_BLC<21> A_BLC<20> A_BLC<23> A_BLC<22> A_BLT<21> A_BLT<20> A_BLT<23> A_BLT<22> A_LWL<191> A_LWL<190> A_LWL<189> A_LWL<188> A_LWL<187> A_LWL<186> A_LWL<185> A_LWL<184> A_LWL<183> A_LWL<182> A_LWL<181> A_LWL<180> A_LWL<179> A_LWL<178> A_LWL<177> A_LWL<176> A_RWL<191> A_RWL<190> A_RWL<189> A_RWL<188> A_RWL<187> A_RWL<186> A_RWL<185> A_RWL<184> A_RWL<183> A_RWL<182> A_RWL<181> A_RWL<180> A_RWL<179> A_RWL<178> A_RWL<177> A_RWL<176> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<11> A_BLC<19> A_BLC<18> A_BLC<21> A_BLC<20> A_BLT<19> A_BLT<18> A_BLT<21> A_BLT<20> A_LWL<175> A_LWL<174> A_LWL<173> A_LWL<172> A_LWL<171> A_LWL<170> A_LWL<169> A_LWL<168> A_LWL<167> A_LWL<166> A_LWL<165> A_LWL<164> A_LWL<163> A_LWL<162> A_LWL<161> A_LWL<160> A_RWL<175> A_RWL<174> A_RWL<173> A_RWL<172> A_RWL<171> A_RWL<170> A_RWL<169> A_RWL<168> A_RWL<167> A_RWL<166> A_RWL<165> A_RWL<164> A_RWL<163> A_RWL<162> A_RWL<161> A_RWL<160> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<10> A_BLC<17> A_BLC<16> A_BLC<19> A_BLC<18> A_BLT<17> A_BLT<16> A_BLT<19> A_BLT<18> A_LWL<159> A_LWL<158> A_LWL<157> A_LWL<156> A_LWL<155> A_LWL<154> A_LWL<153> A_LWL<152> A_LWL<151> A_LWL<150> A_LWL<149> A_LWL<148> A_LWL<147> A_LWL<146> A_LWL<145> A_LWL<144> A_RWL<159> A_RWL<158> A_RWL<157> A_RWL<156> A_RWL<155> A_RWL<154> A_RWL<153> A_RWL<152> A_RWL<151> A_RWL<150> A_RWL<149> A_RWL<148> A_RWL<147> A_RWL<146> A_RWL<145> A_RWL<144> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<9> A_BLC<15> A_BLC<14> A_BLC<17> A_BLC<16> A_BLT<15> A_BLT<14> A_BLT<17> A_BLT<16> A_LWL<143> A_LWL<142> A_LWL<141> A_LWL<140> A_LWL<139> A_LWL<138> A_LWL<137> A_LWL<136> A_LWL<135> A_LWL<134> A_LWL<133> A_LWL<132> A_LWL<131> A_LWL<130> A_LWL<129> A_LWL<128> A_RWL<143> A_RWL<142> A_RWL<141> A_RWL<140> A_RWL<139> A_RWL<138> A_RWL<137> A_RWL<136> A_RWL<135> A_RWL<134> A_RWL<133> A_RWL<132> A_RWL<131> A_RWL<130> A_RWL<129> A_RWL<128> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<8> A_BLC<13> A_BLC<12> A_BLC<15> A_BLC<14> A_BLT<13> A_BLT<12> A_BLT<15> A_BLT<14> A_LWL<127> A_LWL<126> A_LWL<125> A_LWL<124> A_LWL<123> A_LWL<122> A_LWL<121> A_LWL<120> A_LWL<119> A_LWL<118> A_LWL<117> A_LWL<116> A_LWL<115> A_LWL<114> A_LWL<113> A_LWL<112> A_RWL<127> A_RWL<126> A_RWL<125> A_RWL<124> A_RWL<123> A_RWL<122> A_RWL<121> A_RWL<120> A_RWL<119> A_RWL<118> A_RWL<117> A_RWL<116> A_RWL<115> A_RWL<114> A_RWL<113> A_RWL<112> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<7> A_BLC<11> A_BLC<10> A_BLC<13> A_BLC<12> A_BLT<11> A_BLT<10> A_BLT<13> A_BLT<12> A_LWL<111> A_LWL<110> A_LWL<109> A_LWL<108> A_LWL<107> A_LWL<106> A_LWL<105> A_LWL<104> A_LWL<103> A_LWL<102> A_LWL<101> A_LWL<100> A_LWL<99> A_LWL<98> A_LWL<97> A_LWL<96> A_RWL<111> A_RWL<110> A_RWL<109> A_RWL<108> A_RWL<107> A_RWL<106> A_RWL<105> A_RWL<104> A_RWL<103> A_RWL<102> A_RWL<101> A_RWL<100> A_RWL<99> A_RWL<98> A_RWL<97> A_RWL<96> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<6> A_BLC<9> A_BLC<8> A_BLC<11> A_BLC<10> A_BLT<9> A_BLT<8> A_BLT<11> A_BLT<10> A_LWL<95> A_LWL<94> A_LWL<93> A_LWL<92> A_LWL<91> A_LWL<90> A_LWL<89> A_LWL<88> A_LWL<87> A_LWL<86> A_LWL<85> A_LWL<84> A_LWL<83> A_LWL<82> A_LWL<81> A_LWL<80> A_RWL<95> A_RWL<94> A_RWL<93> A_RWL<92> A_RWL<91> A_RWL<90> A_RWL<89> A_RWL<88> A_RWL<87> A_RWL<86> A_RWL<85> A_RWL<84> A_RWL<83> A_RWL<82> A_RWL<81> A_RWL<80> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<5> A_BLC<7> A_BLC<6> A_BLC<9> A_BLC<8> A_BLT<7> A_BLT<6> A_BLT<9> A_BLT<8> A_LWL<79> A_LWL<78> A_LWL<77> A_LWL<76> A_LWL<75> A_LWL<74> A_LWL<73> A_LWL<72> A_LWL<71> A_LWL<70> A_LWL<69> A_LWL<68> A_LWL<67> A_LWL<66> A_LWL<65> A_LWL<64> A_RWL<79> A_RWL<78> A_RWL<77> A_RWL<76> A_RWL<75> A_RWL<74> A_RWL<73> A_RWL<72> A_RWL<71> A_RWL<70> A_RWL<69> A_RWL<68> A_RWL<67> A_RWL<66> A_RWL<65> A_RWL<64> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<4> A_BLC<5> A_BLC<4> A_BLC<7> A_BLC<6> A_BLT<5> A_BLT<4> A_BLT<7> A_BLT<6> A_LWL<63> A_LWL<62> A_LWL<61> A_LWL<60> A_LWL<59> A_LWL<58> A_LWL<57> A_LWL<56> A_LWL<55> A_LWL<54> A_LWL<53> A_LWL<52> A_LWL<51> A_LWL<50> A_LWL<49> A_LWL<48> A_RWL<63> A_RWL<62> A_RWL<61> A_RWL<60> A_RWL<59> A_RWL<58> A_RWL<57> A_RWL<56> A_RWL<55> A_RWL<54> A_RWL<53> A_RWL<52> A_RWL<51> A_RWL<50> A_RWL<49> A_RWL<48> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<3> A_BLC<3> A_BLC<2> A_BLC<5> A_BLC<4> A_BLT<3> A_BLT<2> A_BLT<5> A_BLT<4> A_LWL<47> A_LWL<46> A_LWL<45> A_LWL<44> A_LWL<43> A_LWL<42> A_LWL<41> A_LWL<40> A_LWL<39> A_LWL<38> A_LWL<37> A_LWL<36> A_LWL<35> A_LWL<34> A_LWL<33> A_LWL<32> A_RWL<47> A_RWL<46> A_RWL<45> A_RWL<44> A_RWL<43> A_RWL<42> A_RWL<41> A_RWL<40> A_RWL<39> A_RWL<38> A_RWL<37> A_RWL<36> A_RWL<35> A_RWL<34> A_RWL<33> A_RWL<32> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<2> A_BLC<1> A_BLC<0> A_BLC<3> A_BLC<2> A_BLT<1> A_BLT<0> A_BLT<3> A_BLT<2> A_LWL<31> A_LWL<30> A_LWL<29> A_LWL<28> A_LWL<27> A_LWL<26> A_LWL<25> A_LWL<24> A_LWL<23> A_LWL<22> A_LWL<21> A_LWL<20> A_LWL<19> A_LWL<18> A_LWL<17> A_LWL<16> A_RWL<31> A_RWL<30> A_RWL<29> A_RWL<28> A_RWL<27> A_RWL<26> A_RWL<25> A_RWL<24> A_RWL<23> A_RWL<22> A_RWL<21> A_RWL<20> A_RWL<19> A_RWL<18> A_RWL<17> A_RWL<16> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XRAM<1> A_BLC_BOT<1> A_BLC_BOT<0> A_BLC<1> A_BLC<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT<1> A_BLT<0> A_LWL<15> A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_SRAM
XEDGE<1> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT_TOP<1> A_BLT_TOP<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_TB
XEDGE<0> A_BLC_BOT<1> A_BLC_BOT<0> A_BLT_BOT<1> A_BLT_BOT<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_TB
.ENDS




.SUBCKT RM_IHPSG13_1024x64_c2_1P_MATRIX_pcell_1 A_BLC<127> A_BLC<126> A_BLC<125> A_BLC<124> A_BLC<123> A_BLC<122> A_BLC<121> A_BLC<120> A_BLC<119> A_BLC<118> A_BLC<117> A_BLC<116> A_BLC<115> A_BLC<114> A_BLC<113> A_BLC<112> A_BLC<111> A_BLC<110> A_BLC<109> A_BLC<108> A_BLC<107> A_BLC<106> A_BLC<105> A_BLC<104> A_BLC<103> A_BLC<102> A_BLC<101> A_BLC<100> A_BLC<99> A_BLC<98> A_BLC<97> A_BLC<96> A_BLC<95> A_BLC<94> A_BLC<93> A_BLC<92> A_BLC<91> A_BLC<90> A_BLC<89> A_BLC<88> A_BLC<87> A_BLC<86> A_BLC<85> A_BLC<84> A_BLC<83> A_BLC<82> A_BLC<81> A_BLC<80> A_BLC<79> A_BLC<78> A_BLC<77> A_BLC<76> A_BLC<75> A_BLC<74> A_BLC<73> A_BLC<72> A_BLC<71> A_BLC<70> A_BLC<69> A_BLC<68> A_BLC<67> A_BLC<66> A_BLC<65> A_BLC<64> A_BLC<63> A_BLC<62> A_BLC<61> A_BLC<60> A_BLC<59> A_BLC<58> A_BLC<57> A_BLC<56> A_BLC<55> A_BLC<54> A_BLC<53> A_BLC<52> A_BLC<51> A_BLC<50> A_BLC<49> A_BLC<48> A_BLC<47> A_BLC<46> A_BLC<45> A_BLC<44> A_BLC<43> A_BLC<42> A_BLC<41> A_BLC<40> A_BLC<39> A_BLC<38> A_BLC<37> A_BLC<36> A_BLC<35> A_BLC<34> A_BLC<33> A_BLC<32> A_BLC<31> A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<127> A_BLT<126> A_BLT<125> A_BLT<124> A_BLT<123> A_BLT<122> A_BLT<121> A_BLT<120> A_BLT<119> A_BLT<118> A_BLT<117> A_BLT<116> A_BLT<115> A_BLT<114> A_BLT<113> A_BLT<112> A_BLT<111> A_BLT<110> A_BLT<109> A_BLT<108> A_BLT<107> A_BLT<106> A_BLT<105> A_BLT<104> A_BLT<103> A_BLT<102> A_BLT<101> A_BLT<100> A_BLT<99> A_BLT<98> A_BLT<97> A_BLT<96> A_BLT<95> A_BLT<94> A_BLT<93> A_BLT<92> A_BLT<91> A_BLT<90> A_BLT<89> A_BLT<88> A_BLT<87> A_BLT<86> A_BLT<85> A_BLT<84> A_BLT<83> A_BLT<82> A_BLT<81> A_BLT<80> A_BLT<79> A_BLT<78> A_BLT<77> A_BLT<76> A_BLT<75> A_BLT<74> A_BLT<73> A_BLT<72> A_BLT<71> A_BLT<70> A_BLT<69> A_BLT<68> A_BLT<67> A_BLT<66> A_BLT<65> A_BLT<64> A_BLT<63> A_BLT<62> A_BLT<61> A_BLT<60> A_BLT<59> A_BLT<58> A_BLT<57> A_BLT<56> A_BLT<55> A_BLT<54> A_BLT<53> A_BLT<52> A_BLT<51> A_BLT<50> A_BLT<49> A_BLT<48> A_BLT<47> A_BLT<46> A_BLT<45> A_BLT<44> A_BLT<43> A_BLT<42> A_BLT<41> A_BLT<40> A_BLT<39> A_BLT<38> A_BLT<37> A_BLT<36> A_BLT<35> A_BLT<34> A_BLT<33> A_BLT<32> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_WL<255> A_WL<254> A_WL<253> A_WL<252> A_WL<251> A_WL<250> A_WL<249> A_WL<248> A_WL<247> A_WL<246> A_WL<245> A_WL<244> A_WL<243> A_WL<242> A_WL<241> A_WL<240> A_WL<239> A_WL<238> A_WL<237> A_WL<236> A_WL<235> A_WL<234> A_WL<233> A_WL<232> A_WL<231> A_WL<230> A_WL<229> A_WL<228> A_WL<227> A_WL<226> A_WL<225> A_WL<224> A_WL<223> A_WL<222> A_WL<221> A_WL<220> A_WL<219> A_WL<218> A_WL<217> A_WL<216> A_WL<215> A_WL<214> A_WL<213> A_WL<212> A_WL<211> A_WL<210> A_WL<209> A_WL<208> A_WL<207> A_WL<206> A_WL<205> A_WL<204> A_WL<203> A_WL<202> A_WL<201> A_WL<200> A_WL<199> A_WL<198> A_WL<197> A_WL<196> A_WL<195> A_WL<194> A_WL<193> A_WL<192> A_WL<191> A_WL<190> A_WL<189> A_WL<188> A_WL<187> A_WL<186> A_WL<185> A_WL<184> A_WL<183> A_WL<182> A_WL<181> A_WL<180> A_WL<179> A_WL<178> A_WL<177> A_WL<176> A_WL<175> A_WL<174> A_WL<173> A_WL<172> A_WL<171> A_WL<170> A_WL<169> A_WL<168> A_WL<167> A_WL<166> A_WL<165> A_WL<164> A_WL<163> A_WL<162> A_WL<161> A_WL<160> A_WL<159> A_WL<158> A_WL<157> A_WL<156> A_WL<155> A_WL<154> A_WL<153> A_WL<152> A_WL<151> A_WL<150> A_WL<149> A_WL<148> A_WL<147> A_WL<146> A_WL<145> A_WL<144> A_WL<143> A_WL<142> A_WL<141> A_WL<140> A_WL<139> A_WL<138> A_WL<137> A_WL<136> A_WL<135> A_WL<134> A_WL<133> A_WL<132> A_WL<131> A_WL<130> A_WL<129> A_WL<128> A_WL<127> A_WL<126> A_WL<125> A_WL<124> A_WL<123> A_WL<122> A_WL<121> A_WL<120> A_WL<119> A_WL<118> A_WL<117> A_WL<116> A_WL<115> A_WL<114> A_WL<113> A_WL<112> A_WL<111> A_WL<110> A_WL<109> A_WL<108> A_WL<107> A_WL<106> A_WL<105> A_WL<104> A_WL<103> A_WL<102> A_WL<101> A_WL<100> A_WL<99> A_WL<98> A_WL<97> A_WL<96> A_WL<95> A_WL<94> A_WL<93> A_WL<92> A_WL<91> A_WL<90> A_WL<89> A_WL<88> A_WL<87> A_WL<86> A_WL<85> A_WL<84> A_WL<83> A_WL<82> A_WL<81> A_WL<80> A_WL<79> A_WL<78> A_WL<77> A_WL<76> A_WL<75> A_WL<74> A_WL<73> A_WL<72> A_WL<71> A_WL<70> A_WL<69> A_WL<68> A_WL<67> A_WL<66> A_WL<65> A_WL<64> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS
XCORNER<3> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_CORNER
XCORNER<2> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_CORNER
XCORNER<1> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_CORNER
XCORNER<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_CORNER
XRAMEDGE_L<15> A_WL<255> A_WL<254> A_WL<253> A_WL<252> A_WL<251> A_WL<250> A_WL<249> A_WL<248> A_WL<247> A_WL<246> A_WL<245> A_WL<244> A_WL<243> A_WL<242> A_WL<241> A_WL<240> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<14> A_WL<239> A_WL<238> A_WL<237> A_WL<236> A_WL<235> A_WL<234> A_WL<233> A_WL<232> A_WL<231> A_WL<230> A_WL<229> A_WL<228> A_WL<227> A_WL<226> A_WL<225> A_WL<224> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<13> A_WL<223> A_WL<222> A_WL<221> A_WL<220> A_WL<219> A_WL<218> A_WL<217> A_WL<216> A_WL<215> A_WL<214> A_WL<213> A_WL<212> A_WL<211> A_WL<210> A_WL<209> A_WL<208> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<12> A_WL<207> A_WL<206> A_WL<205> A_WL<204> A_WL<203> A_WL<202> A_WL<201> A_WL<200> A_WL<199> A_WL<198> A_WL<197> A_WL<196> A_WL<195> A_WL<194> A_WL<193> A_WL<192> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<11> A_WL<191> A_WL<190> A_WL<189> A_WL<188> A_WL<187> A_WL<186> A_WL<185> A_WL<184> A_WL<183> A_WL<182> A_WL<181> A_WL<180> A_WL<179> A_WL<178> A_WL<177> A_WL<176> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<10> A_WL<175> A_WL<174> A_WL<173> A_WL<172> A_WL<171> A_WL<170> A_WL<169> A_WL<168> A_WL<167> A_WL<166> A_WL<165> A_WL<164> A_WL<163> A_WL<162> A_WL<161> A_WL<160> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<9> A_WL<159> A_WL<158> A_WL<157> A_WL<156> A_WL<155> A_WL<154> A_WL<153> A_WL<152> A_WL<151> A_WL<150> A_WL<149> A_WL<148> A_WL<147> A_WL<146> A_WL<145> A_WL<144> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<8> A_WL<143> A_WL<142> A_WL<141> A_WL<140> A_WL<139> A_WL<138> A_WL<137> A_WL<136> A_WL<135> A_WL<134> A_WL<133> A_WL<132> A_WL<131> A_WL<130> A_WL<129> A_WL<128> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<7> A_WL<127> A_WL<126> A_WL<125> A_WL<124> A_WL<123> A_WL<122> A_WL<121> A_WL<120> A_WL<119> A_WL<118> A_WL<117> A_WL<116> A_WL<115> A_WL<114> A_WL<113> A_WL<112> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<6> A_WL<111> A_WL<110> A_WL<109> A_WL<108> A_WL<107> A_WL<106> A_WL<105> A_WL<104> A_WL<103> A_WL<102> A_WL<101> A_WL<100> A_WL<99> A_WL<98> A_WL<97> A_WL<96> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<5> A_WL<95> A_WL<94> A_WL<93> A_WL<92> A_WL<91> A_WL<90> A_WL<89> A_WL<88> A_WL<87> A_WL<86> A_WL<85> A_WL<84> A_WL<83> A_WL<82> A_WL<81> A_WL<80> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<4> A_WL<79> A_WL<78> A_WL<77> A_WL<76> A_WL<75> A_WL<74> A_WL<73> A_WL<72> A_WL<71> A_WL<70> A_WL<69> A_WL<68> A_WL<67> A_WL<66> A_WL<65> A_WL<64> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<3> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<2> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<1> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<0> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<15> A_IWL<16383> A_IWL<16382> A_IWL<16381> A_IWL<16380> A_IWL<16379> A_IWL<16378> A_IWL<16377> A_IWL<16376> A_IWL<16375> A_IWL<16374> A_IWL<16373> A_IWL<16372> A_IWL<16371> A_IWL<16370> A_IWL<16369> A_IWL<16368> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<14> A_IWL<16367> A_IWL<16366> A_IWL<16365> A_IWL<16364> A_IWL<16363> A_IWL<16362> A_IWL<16361> A_IWL<16360> A_IWL<16359> A_IWL<16358> A_IWL<16357> A_IWL<16356> A_IWL<16355> A_IWL<16354> A_IWL<16353> A_IWL<16352> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<13> A_IWL<16351> A_IWL<16350> A_IWL<16349> A_IWL<16348> A_IWL<16347> A_IWL<16346> A_IWL<16345> A_IWL<16344> A_IWL<16343> A_IWL<16342> A_IWL<16341> A_IWL<16340> A_IWL<16339> A_IWL<16338> A_IWL<16337> A_IWL<16336> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<12> A_IWL<16335> A_IWL<16334> A_IWL<16333> A_IWL<16332> A_IWL<16331> A_IWL<16330> A_IWL<16329> A_IWL<16328> A_IWL<16327> A_IWL<16326> A_IWL<16325> A_IWL<16324> A_IWL<16323> A_IWL<16322> A_IWL<16321> A_IWL<16320> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<11> A_IWL<16319> A_IWL<16318> A_IWL<16317> A_IWL<16316> A_IWL<16315> A_IWL<16314> A_IWL<16313> A_IWL<16312> A_IWL<16311> A_IWL<16310> A_IWL<16309> A_IWL<16308> A_IWL<16307> A_IWL<16306> A_IWL<16305> A_IWL<16304> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<10> A_IWL<16303> A_IWL<16302> A_IWL<16301> A_IWL<16300> A_IWL<16299> A_IWL<16298> A_IWL<16297> A_IWL<16296> A_IWL<16295> A_IWL<16294> A_IWL<16293> A_IWL<16292> A_IWL<16291> A_IWL<16290> A_IWL<16289> A_IWL<16288> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<9> A_IWL<16287> A_IWL<16286> A_IWL<16285> A_IWL<16284> A_IWL<16283> A_IWL<16282> A_IWL<16281> A_IWL<16280> A_IWL<16279> A_IWL<16278> A_IWL<16277> A_IWL<16276> A_IWL<16275> A_IWL<16274> A_IWL<16273> A_IWL<16272> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<8> A_IWL<16271> A_IWL<16270> A_IWL<16269> A_IWL<16268> A_IWL<16267> A_IWL<16266> A_IWL<16265> A_IWL<16264> A_IWL<16263> A_IWL<16262> A_IWL<16261> A_IWL<16260> A_IWL<16259> A_IWL<16258> A_IWL<16257> A_IWL<16256> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<7> A_IWL<16255> A_IWL<16254> A_IWL<16253> A_IWL<16252> A_IWL<16251> A_IWL<16250> A_IWL<16249> A_IWL<16248> A_IWL<16247> A_IWL<16246> A_IWL<16245> A_IWL<16244> A_IWL<16243> A_IWL<16242> A_IWL<16241> A_IWL<16240> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<6> A_IWL<16239> A_IWL<16238> A_IWL<16237> A_IWL<16236> A_IWL<16235> A_IWL<16234> A_IWL<16233> A_IWL<16232> A_IWL<16231> A_IWL<16230> A_IWL<16229> A_IWL<16228> A_IWL<16227> A_IWL<16226> A_IWL<16225> A_IWL<16224> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<5> A_IWL<16223> A_IWL<16222> A_IWL<16221> A_IWL<16220> A_IWL<16219> A_IWL<16218> A_IWL<16217> A_IWL<16216> A_IWL<16215> A_IWL<16214> A_IWL<16213> A_IWL<16212> A_IWL<16211> A_IWL<16210> A_IWL<16209> A_IWL<16208> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<4> A_IWL<16207> A_IWL<16206> A_IWL<16205> A_IWL<16204> A_IWL<16203> A_IWL<16202> A_IWL<16201> A_IWL<16200> A_IWL<16199> A_IWL<16198> A_IWL<16197> A_IWL<16196> A_IWL<16195> A_IWL<16194> A_IWL<16193> A_IWL<16192> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<3> A_IWL<16191> A_IWL<16190> A_IWL<16189> A_IWL<16188> A_IWL<16187> A_IWL<16186> A_IWL<16185> A_IWL<16184> A_IWL<16183> A_IWL<16182> A_IWL<16181> A_IWL<16180> A_IWL<16179> A_IWL<16178> A_IWL<16177> A_IWL<16176> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<2> A_IWL<16175> A_IWL<16174> A_IWL<16173> A_IWL<16172> A_IWL<16171> A_IWL<16170> A_IWL<16169> A_IWL<16168> A_IWL<16167> A_IWL<16166> A_IWL<16165> A_IWL<16164> A_IWL<16163> A_IWL<16162> A_IWL<16161> A_IWL<16160> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<1> A_IWL<16159> A_IWL<16158> A_IWL<16157> A_IWL<16156> A_IWL<16155> A_IWL<16154> A_IWL<16153> A_IWL<16152> A_IWL<16151> A_IWL<16150> A_IWL<16149> A_IWL<16148> A_IWL<16147> A_IWL<16146> A_IWL<16145> A_IWL<16144> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<0> A_IWL<16143> A_IWL<16142> A_IWL<16141> A_IWL<16140> A_IWL<16139> A_IWL<16138> A_IWL<16137> A_IWL<16136> A_IWL<16135> A_IWL<16134> A_IWL<16133> A_IWL<16132> A_IWL<16131> A_IWL<16130> A_IWL<16129> A_IWL<16128> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_BITKIT_16x2_EDGE_LR
XCOL<63> A_BLC<127> A_BLC<126> A_BLC_TOP<127> A_BLC_TOP<126> A_BLT<127> A_BLT<126> A_BLT_TOP<127> A_BLT_TOP<126> A_IWL<16127> A_IWL<16126> A_IWL<16125> A_IWL<16124> A_IWL<16123> A_IWL<16122> A_IWL<16121> A_IWL<16120> A_IWL<16119> A_IWL<16118> A_IWL<16117> A_IWL<16116> A_IWL<16115> A_IWL<16114> A_IWL<16113> A_IWL<16112> A_IWL<16111> A_IWL<16110> A_IWL<16109> A_IWL<16108> A_IWL<16107> A_IWL<16106> A_IWL<16105> A_IWL<16104> A_IWL<16103> A_IWL<16102> A_IWL<16101> A_IWL<16100> A_IWL<16099> A_IWL<16098> A_IWL<16097> A_IWL<16096> A_IWL<16095> A_IWL<16094> A_IWL<16093> A_IWL<16092> A_IWL<16091> A_IWL<16090> A_IWL<16089> A_IWL<16088> A_IWL<16087> A_IWL<16086> A_IWL<16085> A_IWL<16084> A_IWL<16083> A_IWL<16082> A_IWL<16081> A_IWL<16080> A_IWL<16079> A_IWL<16078> A_IWL<16077> A_IWL<16076> A_IWL<16075> A_IWL<16074> A_IWL<16073> A_IWL<16072> A_IWL<16071> A_IWL<16070> A_IWL<16069> A_IWL<16068> A_IWL<16067> A_IWL<16066> A_IWL<16065> A_IWL<16064> A_IWL<16063> A_IWL<16062> A_IWL<16061> A_IWL<16060> A_IWL<16059> A_IWL<16058> A_IWL<16057> A_IWL<16056> A_IWL<16055> A_IWL<16054> A_IWL<16053> A_IWL<16052> A_IWL<16051> A_IWL<16050> A_IWL<16049> A_IWL<16048> A_IWL<16047> A_IWL<16046> A_IWL<16045> A_IWL<16044> A_IWL<16043> A_IWL<16042> A_IWL<16041> A_IWL<16040> A_IWL<16039> A_IWL<16038> A_IWL<16037> A_IWL<16036> A_IWL<16035> A_IWL<16034> A_IWL<16033> A_IWL<16032> A_IWL<16031> A_IWL<16030> A_IWL<16029> A_IWL<16028> A_IWL<16027> A_IWL<16026> A_IWL<16025> A_IWL<16024> A_IWL<16023> A_IWL<16022> A_IWL<16021> A_IWL<16020> A_IWL<16019> A_IWL<16018> A_IWL<16017> A_IWL<16016> A_IWL<16015> A_IWL<16014> A_IWL<16013> A_IWL<16012> A_IWL<16011> A_IWL<16010> A_IWL<16009> A_IWL<16008> A_IWL<16007> A_IWL<16006> A_IWL<16005> A_IWL<16004> A_IWL<16003> A_IWL<16002> A_IWL<16001> A_IWL<16000> A_IWL<15999> A_IWL<15998> A_IWL<15997> A_IWL<15996> A_IWL<15995> A_IWL<15994> A_IWL<15993> A_IWL<15992> A_IWL<15991> A_IWL<15990> A_IWL<15989> A_IWL<15988> A_IWL<15987> A_IWL<15986> A_IWL<15985> A_IWL<15984> A_IWL<15983> A_IWL<15982> A_IWL<15981> A_IWL<15980> A_IWL<15979> A_IWL<15978> A_IWL<15977> A_IWL<15976> A_IWL<15975> A_IWL<15974> A_IWL<15973> A_IWL<15972> A_IWL<15971> A_IWL<15970> A_IWL<15969> A_IWL<15968> A_IWL<15967> A_IWL<15966> A_IWL<15965> A_IWL<15964> A_IWL<15963> A_IWL<15962> A_IWL<15961> A_IWL<15960> A_IWL<15959> A_IWL<15958> A_IWL<15957> A_IWL<15956> A_IWL<15955> A_IWL<15954> A_IWL<15953> A_IWL<15952> A_IWL<15951> A_IWL<15950> A_IWL<15949> A_IWL<15948> A_IWL<15947> A_IWL<15946> A_IWL<15945> A_IWL<15944> A_IWL<15943> A_IWL<15942> A_IWL<15941> A_IWL<15940> A_IWL<15939> A_IWL<15938> A_IWL<15937> A_IWL<15936> A_IWL<15935> A_IWL<15934> A_IWL<15933> A_IWL<15932> A_IWL<15931> A_IWL<15930> A_IWL<15929> A_IWL<15928> A_IWL<15927> A_IWL<15926> A_IWL<15925> A_IWL<15924> A_IWL<15923> A_IWL<15922> A_IWL<15921> A_IWL<15920> A_IWL<15919> A_IWL<15918> A_IWL<15917> A_IWL<15916> A_IWL<15915> A_IWL<15914> A_IWL<15913> A_IWL<15912> A_IWL<15911> A_IWL<15910> A_IWL<15909> A_IWL<15908> A_IWL<15907> A_IWL<15906> A_IWL<15905> A_IWL<15904> A_IWL<15903> A_IWL<15902> A_IWL<15901> A_IWL<15900> A_IWL<15899> A_IWL<15898> A_IWL<15897> A_IWL<15896> A_IWL<15895> A_IWL<15894> A_IWL<15893> A_IWL<15892> A_IWL<15891> A_IWL<15890> A_IWL<15889> A_IWL<15888> A_IWL<15887> A_IWL<15886> A_IWL<15885> A_IWL<15884> A_IWL<15883> A_IWL<15882> A_IWL<15881> A_IWL<15880> A_IWL<15879> A_IWL<15878> A_IWL<15877> A_IWL<15876> A_IWL<15875> A_IWL<15874> A_IWL<15873> A_IWL<15872> A_IWL<16383> A_IWL<16382> A_IWL<16381> A_IWL<16380> A_IWL<16379> A_IWL<16378> A_IWL<16377> A_IWL<16376> A_IWL<16375> A_IWL<16374> A_IWL<16373> A_IWL<16372> A_IWL<16371> A_IWL<16370> A_IWL<16369> A_IWL<16368> A_IWL<16367> A_IWL<16366> A_IWL<16365> A_IWL<16364> A_IWL<16363> A_IWL<16362> A_IWL<16361> A_IWL<16360> A_IWL<16359> A_IWL<16358> A_IWL<16357> A_IWL<16356> A_IWL<16355> A_IWL<16354> A_IWL<16353> A_IWL<16352> A_IWL<16351> A_IWL<16350> A_IWL<16349> A_IWL<16348> A_IWL<16347> A_IWL<16346> A_IWL<16345> A_IWL<16344> A_IWL<16343> A_IWL<16342> A_IWL<16341> A_IWL<16340> A_IWL<16339> A_IWL<16338> A_IWL<16337> A_IWL<16336> A_IWL<16335> A_IWL<16334> A_IWL<16333> A_IWL<16332> A_IWL<16331> A_IWL<16330> A_IWL<16329> A_IWL<16328> A_IWL<16327> A_IWL<16326> A_IWL<16325> A_IWL<16324> A_IWL<16323> A_IWL<16322> A_IWL<16321> A_IWL<16320> A_IWL<16319> A_IWL<16318> A_IWL<16317> A_IWL<16316> A_IWL<16315> A_IWL<16314> A_IWL<16313> A_IWL<16312> A_IWL<16311> A_IWL<16310> A_IWL<16309> A_IWL<16308> A_IWL<16307> A_IWL<16306> A_IWL<16305> A_IWL<16304> A_IWL<16303> A_IWL<16302> A_IWL<16301> A_IWL<16300> A_IWL<16299> A_IWL<16298> A_IWL<16297> A_IWL<16296> A_IWL<16295> A_IWL<16294> A_IWL<16293> A_IWL<16292> A_IWL<16291> A_IWL<16290> A_IWL<16289> A_IWL<16288> A_IWL<16287> A_IWL<16286> A_IWL<16285> A_IWL<16284> A_IWL<16283> A_IWL<16282> A_IWL<16281> A_IWL<16280> A_IWL<16279> A_IWL<16278> A_IWL<16277> A_IWL<16276> A_IWL<16275> A_IWL<16274> A_IWL<16273> A_IWL<16272> A_IWL<16271> A_IWL<16270> A_IWL<16269> A_IWL<16268> A_IWL<16267> A_IWL<16266> A_IWL<16265> A_IWL<16264> A_IWL<16263> A_IWL<16262> A_IWL<16261> A_IWL<16260> A_IWL<16259> A_IWL<16258> A_IWL<16257> A_IWL<16256> A_IWL<16255> A_IWL<16254> A_IWL<16253> A_IWL<16252> A_IWL<16251> A_IWL<16250> A_IWL<16249> A_IWL<16248> A_IWL<16247> A_IWL<16246> A_IWL<16245> A_IWL<16244> A_IWL<16243> A_IWL<16242> A_IWL<16241> A_IWL<16240> A_IWL<16239> A_IWL<16238> A_IWL<16237> A_IWL<16236> A_IWL<16235> A_IWL<16234> A_IWL<16233> A_IWL<16232> A_IWL<16231> A_IWL<16230> A_IWL<16229> A_IWL<16228> A_IWL<16227> A_IWL<16226> A_IWL<16225> A_IWL<16224> A_IWL<16223> A_IWL<16222> A_IWL<16221> A_IWL<16220> A_IWL<16219> A_IWL<16218> A_IWL<16217> A_IWL<16216> A_IWL<16215> A_IWL<16214> A_IWL<16213> A_IWL<16212> A_IWL<16211> A_IWL<16210> A_IWL<16209> A_IWL<16208> A_IWL<16207> A_IWL<16206> A_IWL<16205> A_IWL<16204> A_IWL<16203> A_IWL<16202> A_IWL<16201> A_IWL<16200> A_IWL<16199> A_IWL<16198> A_IWL<16197> A_IWL<16196> A_IWL<16195> A_IWL<16194> A_IWL<16193> A_IWL<16192> A_IWL<16191> A_IWL<16190> A_IWL<16189> A_IWL<16188> A_IWL<16187> A_IWL<16186> A_IWL<16185> A_IWL<16184> A_IWL<16183> A_IWL<16182> A_IWL<16181> A_IWL<16180> A_IWL<16179> A_IWL<16178> A_IWL<16177> A_IWL<16176> A_IWL<16175> A_IWL<16174> A_IWL<16173> A_IWL<16172> A_IWL<16171> A_IWL<16170> A_IWL<16169> A_IWL<16168> A_IWL<16167> A_IWL<16166> A_IWL<16165> A_IWL<16164> A_IWL<16163> A_IWL<16162> A_IWL<16161> A_IWL<16160> A_IWL<16159> A_IWL<16158> A_IWL<16157> A_IWL<16156> A_IWL<16155> A_IWL<16154> A_IWL<16153> A_IWL<16152> A_IWL<16151> A_IWL<16150> A_IWL<16149> A_IWL<16148> A_IWL<16147> A_IWL<16146> A_IWL<16145> A_IWL<16144> A_IWL<16143> A_IWL<16142> A_IWL<16141> A_IWL<16140> A_IWL<16139> A_IWL<16138> A_IWL<16137> A_IWL<16136> A_IWL<16135> A_IWL<16134> A_IWL<16133> A_IWL<16132> A_IWL<16131> A_IWL<16130> A_IWL<16129> A_IWL<16128> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<62> A_BLC<125> A_BLC<124> A_BLC_TOP<125> A_BLC_TOP<124> A_BLT<125> A_BLT<124> A_BLT_TOP<125> A_BLT_TOP<124> A_IWL<15871> A_IWL<15870> A_IWL<15869> A_IWL<15868> A_IWL<15867> A_IWL<15866> A_IWL<15865> A_IWL<15864> A_IWL<15863> A_IWL<15862> A_IWL<15861> A_IWL<15860> A_IWL<15859> A_IWL<15858> A_IWL<15857> A_IWL<15856> A_IWL<15855> A_IWL<15854> A_IWL<15853> A_IWL<15852> A_IWL<15851> A_IWL<15850> A_IWL<15849> A_IWL<15848> A_IWL<15847> A_IWL<15846> A_IWL<15845> A_IWL<15844> A_IWL<15843> A_IWL<15842> A_IWL<15841> A_IWL<15840> A_IWL<15839> A_IWL<15838> A_IWL<15837> A_IWL<15836> A_IWL<15835> A_IWL<15834> A_IWL<15833> A_IWL<15832> A_IWL<15831> A_IWL<15830> A_IWL<15829> A_IWL<15828> A_IWL<15827> A_IWL<15826> A_IWL<15825> A_IWL<15824> A_IWL<15823> A_IWL<15822> A_IWL<15821> A_IWL<15820> A_IWL<15819> A_IWL<15818> A_IWL<15817> A_IWL<15816> A_IWL<15815> A_IWL<15814> A_IWL<15813> A_IWL<15812> A_IWL<15811> A_IWL<15810> A_IWL<15809> A_IWL<15808> A_IWL<15807> A_IWL<15806> A_IWL<15805> A_IWL<15804> A_IWL<15803> A_IWL<15802> A_IWL<15801> A_IWL<15800> A_IWL<15799> A_IWL<15798> A_IWL<15797> A_IWL<15796> A_IWL<15795> A_IWL<15794> A_IWL<15793> A_IWL<15792> A_IWL<15791> A_IWL<15790> A_IWL<15789> A_IWL<15788> A_IWL<15787> A_IWL<15786> A_IWL<15785> A_IWL<15784> A_IWL<15783> A_IWL<15782> A_IWL<15781> A_IWL<15780> A_IWL<15779> A_IWL<15778> A_IWL<15777> A_IWL<15776> A_IWL<15775> A_IWL<15774> A_IWL<15773> A_IWL<15772> A_IWL<15771> A_IWL<15770> A_IWL<15769> A_IWL<15768> A_IWL<15767> A_IWL<15766> A_IWL<15765> A_IWL<15764> A_IWL<15763> A_IWL<15762> A_IWL<15761> A_IWL<15760> A_IWL<15759> A_IWL<15758> A_IWL<15757> A_IWL<15756> A_IWL<15755> A_IWL<15754> A_IWL<15753> A_IWL<15752> A_IWL<15751> A_IWL<15750> A_IWL<15749> A_IWL<15748> A_IWL<15747> A_IWL<15746> A_IWL<15745> A_IWL<15744> A_IWL<15743> A_IWL<15742> A_IWL<15741> A_IWL<15740> A_IWL<15739> A_IWL<15738> A_IWL<15737> A_IWL<15736> A_IWL<15735> A_IWL<15734> A_IWL<15733> A_IWL<15732> A_IWL<15731> A_IWL<15730> A_IWL<15729> A_IWL<15728> A_IWL<15727> A_IWL<15726> A_IWL<15725> A_IWL<15724> A_IWL<15723> A_IWL<15722> A_IWL<15721> A_IWL<15720> A_IWL<15719> A_IWL<15718> A_IWL<15717> A_IWL<15716> A_IWL<15715> A_IWL<15714> A_IWL<15713> A_IWL<15712> A_IWL<15711> A_IWL<15710> A_IWL<15709> A_IWL<15708> A_IWL<15707> A_IWL<15706> A_IWL<15705> A_IWL<15704> A_IWL<15703> A_IWL<15702> A_IWL<15701> A_IWL<15700> A_IWL<15699> A_IWL<15698> A_IWL<15697> A_IWL<15696> A_IWL<15695> A_IWL<15694> A_IWL<15693> A_IWL<15692> A_IWL<15691> A_IWL<15690> A_IWL<15689> A_IWL<15688> A_IWL<15687> A_IWL<15686> A_IWL<15685> A_IWL<15684> A_IWL<15683> A_IWL<15682> A_IWL<15681> A_IWL<15680> A_IWL<15679> A_IWL<15678> A_IWL<15677> A_IWL<15676> A_IWL<15675> A_IWL<15674> A_IWL<15673> A_IWL<15672> A_IWL<15671> A_IWL<15670> A_IWL<15669> A_IWL<15668> A_IWL<15667> A_IWL<15666> A_IWL<15665> A_IWL<15664> A_IWL<15663> A_IWL<15662> A_IWL<15661> A_IWL<15660> A_IWL<15659> A_IWL<15658> A_IWL<15657> A_IWL<15656> A_IWL<15655> A_IWL<15654> A_IWL<15653> A_IWL<15652> A_IWL<15651> A_IWL<15650> A_IWL<15649> A_IWL<15648> A_IWL<15647> A_IWL<15646> A_IWL<15645> A_IWL<15644> A_IWL<15643> A_IWL<15642> A_IWL<15641> A_IWL<15640> A_IWL<15639> A_IWL<15638> A_IWL<15637> A_IWL<15636> A_IWL<15635> A_IWL<15634> A_IWL<15633> A_IWL<15632> A_IWL<15631> A_IWL<15630> A_IWL<15629> A_IWL<15628> A_IWL<15627> A_IWL<15626> A_IWL<15625> A_IWL<15624> A_IWL<15623> A_IWL<15622> A_IWL<15621> A_IWL<15620> A_IWL<15619> A_IWL<15618> A_IWL<15617> A_IWL<15616> A_IWL<16127> A_IWL<16126> A_IWL<16125> A_IWL<16124> A_IWL<16123> A_IWL<16122> A_IWL<16121> A_IWL<16120> A_IWL<16119> A_IWL<16118> A_IWL<16117> A_IWL<16116> A_IWL<16115> A_IWL<16114> A_IWL<16113> A_IWL<16112> A_IWL<16111> A_IWL<16110> A_IWL<16109> A_IWL<16108> A_IWL<16107> A_IWL<16106> A_IWL<16105> A_IWL<16104> A_IWL<16103> A_IWL<16102> A_IWL<16101> A_IWL<16100> A_IWL<16099> A_IWL<16098> A_IWL<16097> A_IWL<16096> A_IWL<16095> A_IWL<16094> A_IWL<16093> A_IWL<16092> A_IWL<16091> A_IWL<16090> A_IWL<16089> A_IWL<16088> A_IWL<16087> A_IWL<16086> A_IWL<16085> A_IWL<16084> A_IWL<16083> A_IWL<16082> A_IWL<16081> A_IWL<16080> A_IWL<16079> A_IWL<16078> A_IWL<16077> A_IWL<16076> A_IWL<16075> A_IWL<16074> A_IWL<16073> A_IWL<16072> A_IWL<16071> A_IWL<16070> A_IWL<16069> A_IWL<16068> A_IWL<16067> A_IWL<16066> A_IWL<16065> A_IWL<16064> A_IWL<16063> A_IWL<16062> A_IWL<16061> A_IWL<16060> A_IWL<16059> A_IWL<16058> A_IWL<16057> A_IWL<16056> A_IWL<16055> A_IWL<16054> A_IWL<16053> A_IWL<16052> A_IWL<16051> A_IWL<16050> A_IWL<16049> A_IWL<16048> A_IWL<16047> A_IWL<16046> A_IWL<16045> A_IWL<16044> A_IWL<16043> A_IWL<16042> A_IWL<16041> A_IWL<16040> A_IWL<16039> A_IWL<16038> A_IWL<16037> A_IWL<16036> A_IWL<16035> A_IWL<16034> A_IWL<16033> A_IWL<16032> A_IWL<16031> A_IWL<16030> A_IWL<16029> A_IWL<16028> A_IWL<16027> A_IWL<16026> A_IWL<16025> A_IWL<16024> A_IWL<16023> A_IWL<16022> A_IWL<16021> A_IWL<16020> A_IWL<16019> A_IWL<16018> A_IWL<16017> A_IWL<16016> A_IWL<16015> A_IWL<16014> A_IWL<16013> A_IWL<16012> A_IWL<16011> A_IWL<16010> A_IWL<16009> A_IWL<16008> A_IWL<16007> A_IWL<16006> A_IWL<16005> A_IWL<16004> A_IWL<16003> A_IWL<16002> A_IWL<16001> A_IWL<16000> A_IWL<15999> A_IWL<15998> A_IWL<15997> A_IWL<15996> A_IWL<15995> A_IWL<15994> A_IWL<15993> A_IWL<15992> A_IWL<15991> A_IWL<15990> A_IWL<15989> A_IWL<15988> A_IWL<15987> A_IWL<15986> A_IWL<15985> A_IWL<15984> A_IWL<15983> A_IWL<15982> A_IWL<15981> A_IWL<15980> A_IWL<15979> A_IWL<15978> A_IWL<15977> A_IWL<15976> A_IWL<15975> A_IWL<15974> A_IWL<15973> A_IWL<15972> A_IWL<15971> A_IWL<15970> A_IWL<15969> A_IWL<15968> A_IWL<15967> A_IWL<15966> A_IWL<15965> A_IWL<15964> A_IWL<15963> A_IWL<15962> A_IWL<15961> A_IWL<15960> A_IWL<15959> A_IWL<15958> A_IWL<15957> A_IWL<15956> A_IWL<15955> A_IWL<15954> A_IWL<15953> A_IWL<15952> A_IWL<15951> A_IWL<15950> A_IWL<15949> A_IWL<15948> A_IWL<15947> A_IWL<15946> A_IWL<15945> A_IWL<15944> A_IWL<15943> A_IWL<15942> A_IWL<15941> A_IWL<15940> A_IWL<15939> A_IWL<15938> A_IWL<15937> A_IWL<15936> A_IWL<15935> A_IWL<15934> A_IWL<15933> A_IWL<15932> A_IWL<15931> A_IWL<15930> A_IWL<15929> A_IWL<15928> A_IWL<15927> A_IWL<15926> A_IWL<15925> A_IWL<15924> A_IWL<15923> A_IWL<15922> A_IWL<15921> A_IWL<15920> A_IWL<15919> A_IWL<15918> A_IWL<15917> A_IWL<15916> A_IWL<15915> A_IWL<15914> A_IWL<15913> A_IWL<15912> A_IWL<15911> A_IWL<15910> A_IWL<15909> A_IWL<15908> A_IWL<15907> A_IWL<15906> A_IWL<15905> A_IWL<15904> A_IWL<15903> A_IWL<15902> A_IWL<15901> A_IWL<15900> A_IWL<15899> A_IWL<15898> A_IWL<15897> A_IWL<15896> A_IWL<15895> A_IWL<15894> A_IWL<15893> A_IWL<15892> A_IWL<15891> A_IWL<15890> A_IWL<15889> A_IWL<15888> A_IWL<15887> A_IWL<15886> A_IWL<15885> A_IWL<15884> A_IWL<15883> A_IWL<15882> A_IWL<15881> A_IWL<15880> A_IWL<15879> A_IWL<15878> A_IWL<15877> A_IWL<15876> A_IWL<15875> A_IWL<15874> A_IWL<15873> A_IWL<15872> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<61> A_BLC<123> A_BLC<122> A_BLC_TOP<123> A_BLC_TOP<122> A_BLT<123> A_BLT<122> A_BLT_TOP<123> A_BLT_TOP<122> A_IWL<15615> A_IWL<15614> A_IWL<15613> A_IWL<15612> A_IWL<15611> A_IWL<15610> A_IWL<15609> A_IWL<15608> A_IWL<15607> A_IWL<15606> A_IWL<15605> A_IWL<15604> A_IWL<15603> A_IWL<15602> A_IWL<15601> A_IWL<15600> A_IWL<15599> A_IWL<15598> A_IWL<15597> A_IWL<15596> A_IWL<15595> A_IWL<15594> A_IWL<15593> A_IWL<15592> A_IWL<15591> A_IWL<15590> A_IWL<15589> A_IWL<15588> A_IWL<15587> A_IWL<15586> A_IWL<15585> A_IWL<15584> A_IWL<15583> A_IWL<15582> A_IWL<15581> A_IWL<15580> A_IWL<15579> A_IWL<15578> A_IWL<15577> A_IWL<15576> A_IWL<15575> A_IWL<15574> A_IWL<15573> A_IWL<15572> A_IWL<15571> A_IWL<15570> A_IWL<15569> A_IWL<15568> A_IWL<15567> A_IWL<15566> A_IWL<15565> A_IWL<15564> A_IWL<15563> A_IWL<15562> A_IWL<15561> A_IWL<15560> A_IWL<15559> A_IWL<15558> A_IWL<15557> A_IWL<15556> A_IWL<15555> A_IWL<15554> A_IWL<15553> A_IWL<15552> A_IWL<15551> A_IWL<15550> A_IWL<15549> A_IWL<15548> A_IWL<15547> A_IWL<15546> A_IWL<15545> A_IWL<15544> A_IWL<15543> A_IWL<15542> A_IWL<15541> A_IWL<15540> A_IWL<15539> A_IWL<15538> A_IWL<15537> A_IWL<15536> A_IWL<15535> A_IWL<15534> A_IWL<15533> A_IWL<15532> A_IWL<15531> A_IWL<15530> A_IWL<15529> A_IWL<15528> A_IWL<15527> A_IWL<15526> A_IWL<15525> A_IWL<15524> A_IWL<15523> A_IWL<15522> A_IWL<15521> A_IWL<15520> A_IWL<15519> A_IWL<15518> A_IWL<15517> A_IWL<15516> A_IWL<15515> A_IWL<15514> A_IWL<15513> A_IWL<15512> A_IWL<15511> A_IWL<15510> A_IWL<15509> A_IWL<15508> A_IWL<15507> A_IWL<15506> A_IWL<15505> A_IWL<15504> A_IWL<15503> A_IWL<15502> A_IWL<15501> A_IWL<15500> A_IWL<15499> A_IWL<15498> A_IWL<15497> A_IWL<15496> A_IWL<15495> A_IWL<15494> A_IWL<15493> A_IWL<15492> A_IWL<15491> A_IWL<15490> A_IWL<15489> A_IWL<15488> A_IWL<15487> A_IWL<15486> A_IWL<15485> A_IWL<15484> A_IWL<15483> A_IWL<15482> A_IWL<15481> A_IWL<15480> A_IWL<15479> A_IWL<15478> A_IWL<15477> A_IWL<15476> A_IWL<15475> A_IWL<15474> A_IWL<15473> A_IWL<15472> A_IWL<15471> A_IWL<15470> A_IWL<15469> A_IWL<15468> A_IWL<15467> A_IWL<15466> A_IWL<15465> A_IWL<15464> A_IWL<15463> A_IWL<15462> A_IWL<15461> A_IWL<15460> A_IWL<15459> A_IWL<15458> A_IWL<15457> A_IWL<15456> A_IWL<15455> A_IWL<15454> A_IWL<15453> A_IWL<15452> A_IWL<15451> A_IWL<15450> A_IWL<15449> A_IWL<15448> A_IWL<15447> A_IWL<15446> A_IWL<15445> A_IWL<15444> A_IWL<15443> A_IWL<15442> A_IWL<15441> A_IWL<15440> A_IWL<15439> A_IWL<15438> A_IWL<15437> A_IWL<15436> A_IWL<15435> A_IWL<15434> A_IWL<15433> A_IWL<15432> A_IWL<15431> A_IWL<15430> A_IWL<15429> A_IWL<15428> A_IWL<15427> A_IWL<15426> A_IWL<15425> A_IWL<15424> A_IWL<15423> A_IWL<15422> A_IWL<15421> A_IWL<15420> A_IWL<15419> A_IWL<15418> A_IWL<15417> A_IWL<15416> A_IWL<15415> A_IWL<15414> A_IWL<15413> A_IWL<15412> A_IWL<15411> A_IWL<15410> A_IWL<15409> A_IWL<15408> A_IWL<15407> A_IWL<15406> A_IWL<15405> A_IWL<15404> A_IWL<15403> A_IWL<15402> A_IWL<15401> A_IWL<15400> A_IWL<15399> A_IWL<15398> A_IWL<15397> A_IWL<15396> A_IWL<15395> A_IWL<15394> A_IWL<15393> A_IWL<15392> A_IWL<15391> A_IWL<15390> A_IWL<15389> A_IWL<15388> A_IWL<15387> A_IWL<15386> A_IWL<15385> A_IWL<15384> A_IWL<15383> A_IWL<15382> A_IWL<15381> A_IWL<15380> A_IWL<15379> A_IWL<15378> A_IWL<15377> A_IWL<15376> A_IWL<15375> A_IWL<15374> A_IWL<15373> A_IWL<15372> A_IWL<15371> A_IWL<15370> A_IWL<15369> A_IWL<15368> A_IWL<15367> A_IWL<15366> A_IWL<15365> A_IWL<15364> A_IWL<15363> A_IWL<15362> A_IWL<15361> A_IWL<15360> A_IWL<15871> A_IWL<15870> A_IWL<15869> A_IWL<15868> A_IWL<15867> A_IWL<15866> A_IWL<15865> A_IWL<15864> A_IWL<15863> A_IWL<15862> A_IWL<15861> A_IWL<15860> A_IWL<15859> A_IWL<15858> A_IWL<15857> A_IWL<15856> A_IWL<15855> A_IWL<15854> A_IWL<15853> A_IWL<15852> A_IWL<15851> A_IWL<15850> A_IWL<15849> A_IWL<15848> A_IWL<15847> A_IWL<15846> A_IWL<15845> A_IWL<15844> A_IWL<15843> A_IWL<15842> A_IWL<15841> A_IWL<15840> A_IWL<15839> A_IWL<15838> A_IWL<15837> A_IWL<15836> A_IWL<15835> A_IWL<15834> A_IWL<15833> A_IWL<15832> A_IWL<15831> A_IWL<15830> A_IWL<15829> A_IWL<15828> A_IWL<15827> A_IWL<15826> A_IWL<15825> A_IWL<15824> A_IWL<15823> A_IWL<15822> A_IWL<15821> A_IWL<15820> A_IWL<15819> A_IWL<15818> A_IWL<15817> A_IWL<15816> A_IWL<15815> A_IWL<15814> A_IWL<15813> A_IWL<15812> A_IWL<15811> A_IWL<15810> A_IWL<15809> A_IWL<15808> A_IWL<15807> A_IWL<15806> A_IWL<15805> A_IWL<15804> A_IWL<15803> A_IWL<15802> A_IWL<15801> A_IWL<15800> A_IWL<15799> A_IWL<15798> A_IWL<15797> A_IWL<15796> A_IWL<15795> A_IWL<15794> A_IWL<15793> A_IWL<15792> A_IWL<15791> A_IWL<15790> A_IWL<15789> A_IWL<15788> A_IWL<15787> A_IWL<15786> A_IWL<15785> A_IWL<15784> A_IWL<15783> A_IWL<15782> A_IWL<15781> A_IWL<15780> A_IWL<15779> A_IWL<15778> A_IWL<15777> A_IWL<15776> A_IWL<15775> A_IWL<15774> A_IWL<15773> A_IWL<15772> A_IWL<15771> A_IWL<15770> A_IWL<15769> A_IWL<15768> A_IWL<15767> A_IWL<15766> A_IWL<15765> A_IWL<15764> A_IWL<15763> A_IWL<15762> A_IWL<15761> A_IWL<15760> A_IWL<15759> A_IWL<15758> A_IWL<15757> A_IWL<15756> A_IWL<15755> A_IWL<15754> A_IWL<15753> A_IWL<15752> A_IWL<15751> A_IWL<15750> A_IWL<15749> A_IWL<15748> A_IWL<15747> A_IWL<15746> A_IWL<15745> A_IWL<15744> A_IWL<15743> A_IWL<15742> A_IWL<15741> A_IWL<15740> A_IWL<15739> A_IWL<15738> A_IWL<15737> A_IWL<15736> A_IWL<15735> A_IWL<15734> A_IWL<15733> A_IWL<15732> A_IWL<15731> A_IWL<15730> A_IWL<15729> A_IWL<15728> A_IWL<15727> A_IWL<15726> A_IWL<15725> A_IWL<15724> A_IWL<15723> A_IWL<15722> A_IWL<15721> A_IWL<15720> A_IWL<15719> A_IWL<15718> A_IWL<15717> A_IWL<15716> A_IWL<15715> A_IWL<15714> A_IWL<15713> A_IWL<15712> A_IWL<15711> A_IWL<15710> A_IWL<15709> A_IWL<15708> A_IWL<15707> A_IWL<15706> A_IWL<15705> A_IWL<15704> A_IWL<15703> A_IWL<15702> A_IWL<15701> A_IWL<15700> A_IWL<15699> A_IWL<15698> A_IWL<15697> A_IWL<15696> A_IWL<15695> A_IWL<15694> A_IWL<15693> A_IWL<15692> A_IWL<15691> A_IWL<15690> A_IWL<15689> A_IWL<15688> A_IWL<15687> A_IWL<15686> A_IWL<15685> A_IWL<15684> A_IWL<15683> A_IWL<15682> A_IWL<15681> A_IWL<15680> A_IWL<15679> A_IWL<15678> A_IWL<15677> A_IWL<15676> A_IWL<15675> A_IWL<15674> A_IWL<15673> A_IWL<15672> A_IWL<15671> A_IWL<15670> A_IWL<15669> A_IWL<15668> A_IWL<15667> A_IWL<15666> A_IWL<15665> A_IWL<15664> A_IWL<15663> A_IWL<15662> A_IWL<15661> A_IWL<15660> A_IWL<15659> A_IWL<15658> A_IWL<15657> A_IWL<15656> A_IWL<15655> A_IWL<15654> A_IWL<15653> A_IWL<15652> A_IWL<15651> A_IWL<15650> A_IWL<15649> A_IWL<15648> A_IWL<15647> A_IWL<15646> A_IWL<15645> A_IWL<15644> A_IWL<15643> A_IWL<15642> A_IWL<15641> A_IWL<15640> A_IWL<15639> A_IWL<15638> A_IWL<15637> A_IWL<15636> A_IWL<15635> A_IWL<15634> A_IWL<15633> A_IWL<15632> A_IWL<15631> A_IWL<15630> A_IWL<15629> A_IWL<15628> A_IWL<15627> A_IWL<15626> A_IWL<15625> A_IWL<15624> A_IWL<15623> A_IWL<15622> A_IWL<15621> A_IWL<15620> A_IWL<15619> A_IWL<15618> A_IWL<15617> A_IWL<15616> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<60> A_BLC<121> A_BLC<120> A_BLC_TOP<121> A_BLC_TOP<120> A_BLT<121> A_BLT<120> A_BLT_TOP<121> A_BLT_TOP<120> A_IWL<15359> A_IWL<15358> A_IWL<15357> A_IWL<15356> A_IWL<15355> A_IWL<15354> A_IWL<15353> A_IWL<15352> A_IWL<15351> A_IWL<15350> A_IWL<15349> A_IWL<15348> A_IWL<15347> A_IWL<15346> A_IWL<15345> A_IWL<15344> A_IWL<15343> A_IWL<15342> A_IWL<15341> A_IWL<15340> A_IWL<15339> A_IWL<15338> A_IWL<15337> A_IWL<15336> A_IWL<15335> A_IWL<15334> A_IWL<15333> A_IWL<15332> A_IWL<15331> A_IWL<15330> A_IWL<15329> A_IWL<15328> A_IWL<15327> A_IWL<15326> A_IWL<15325> A_IWL<15324> A_IWL<15323> A_IWL<15322> A_IWL<15321> A_IWL<15320> A_IWL<15319> A_IWL<15318> A_IWL<15317> A_IWL<15316> A_IWL<15315> A_IWL<15314> A_IWL<15313> A_IWL<15312> A_IWL<15311> A_IWL<15310> A_IWL<15309> A_IWL<15308> A_IWL<15307> A_IWL<15306> A_IWL<15305> A_IWL<15304> A_IWL<15303> A_IWL<15302> A_IWL<15301> A_IWL<15300> A_IWL<15299> A_IWL<15298> A_IWL<15297> A_IWL<15296> A_IWL<15295> A_IWL<15294> A_IWL<15293> A_IWL<15292> A_IWL<15291> A_IWL<15290> A_IWL<15289> A_IWL<15288> A_IWL<15287> A_IWL<15286> A_IWL<15285> A_IWL<15284> A_IWL<15283> A_IWL<15282> A_IWL<15281> A_IWL<15280> A_IWL<15279> A_IWL<15278> A_IWL<15277> A_IWL<15276> A_IWL<15275> A_IWL<15274> A_IWL<15273> A_IWL<15272> A_IWL<15271> A_IWL<15270> A_IWL<15269> A_IWL<15268> A_IWL<15267> A_IWL<15266> A_IWL<15265> A_IWL<15264> A_IWL<15263> A_IWL<15262> A_IWL<15261> A_IWL<15260> A_IWL<15259> A_IWL<15258> A_IWL<15257> A_IWL<15256> A_IWL<15255> A_IWL<15254> A_IWL<15253> A_IWL<15252> A_IWL<15251> A_IWL<15250> A_IWL<15249> A_IWL<15248> A_IWL<15247> A_IWL<15246> A_IWL<15245> A_IWL<15244> A_IWL<15243> A_IWL<15242> A_IWL<15241> A_IWL<15240> A_IWL<15239> A_IWL<15238> A_IWL<15237> A_IWL<15236> A_IWL<15235> A_IWL<15234> A_IWL<15233> A_IWL<15232> A_IWL<15231> A_IWL<15230> A_IWL<15229> A_IWL<15228> A_IWL<15227> A_IWL<15226> A_IWL<15225> A_IWL<15224> A_IWL<15223> A_IWL<15222> A_IWL<15221> A_IWL<15220> A_IWL<15219> A_IWL<15218> A_IWL<15217> A_IWL<15216> A_IWL<15215> A_IWL<15214> A_IWL<15213> A_IWL<15212> A_IWL<15211> A_IWL<15210> A_IWL<15209> A_IWL<15208> A_IWL<15207> A_IWL<15206> A_IWL<15205> A_IWL<15204> A_IWL<15203> A_IWL<15202> A_IWL<15201> A_IWL<15200> A_IWL<15199> A_IWL<15198> A_IWL<15197> A_IWL<15196> A_IWL<15195> A_IWL<15194> A_IWL<15193> A_IWL<15192> A_IWL<15191> A_IWL<15190> A_IWL<15189> A_IWL<15188> A_IWL<15187> A_IWL<15186> A_IWL<15185> A_IWL<15184> A_IWL<15183> A_IWL<15182> A_IWL<15181> A_IWL<15180> A_IWL<15179> A_IWL<15178> A_IWL<15177> A_IWL<15176> A_IWL<15175> A_IWL<15174> A_IWL<15173> A_IWL<15172> A_IWL<15171> A_IWL<15170> A_IWL<15169> A_IWL<15168> A_IWL<15167> A_IWL<15166> A_IWL<15165> A_IWL<15164> A_IWL<15163> A_IWL<15162> A_IWL<15161> A_IWL<15160> A_IWL<15159> A_IWL<15158> A_IWL<15157> A_IWL<15156> A_IWL<15155> A_IWL<15154> A_IWL<15153> A_IWL<15152> A_IWL<15151> A_IWL<15150> A_IWL<15149> A_IWL<15148> A_IWL<15147> A_IWL<15146> A_IWL<15145> A_IWL<15144> A_IWL<15143> A_IWL<15142> A_IWL<15141> A_IWL<15140> A_IWL<15139> A_IWL<15138> A_IWL<15137> A_IWL<15136> A_IWL<15135> A_IWL<15134> A_IWL<15133> A_IWL<15132> A_IWL<15131> A_IWL<15130> A_IWL<15129> A_IWL<15128> A_IWL<15127> A_IWL<15126> A_IWL<15125> A_IWL<15124> A_IWL<15123> A_IWL<15122> A_IWL<15121> A_IWL<15120> A_IWL<15119> A_IWL<15118> A_IWL<15117> A_IWL<15116> A_IWL<15115> A_IWL<15114> A_IWL<15113> A_IWL<15112> A_IWL<15111> A_IWL<15110> A_IWL<15109> A_IWL<15108> A_IWL<15107> A_IWL<15106> A_IWL<15105> A_IWL<15104> A_IWL<15615> A_IWL<15614> A_IWL<15613> A_IWL<15612> A_IWL<15611> A_IWL<15610> A_IWL<15609> A_IWL<15608> A_IWL<15607> A_IWL<15606> A_IWL<15605> A_IWL<15604> A_IWL<15603> A_IWL<15602> A_IWL<15601> A_IWL<15600> A_IWL<15599> A_IWL<15598> A_IWL<15597> A_IWL<15596> A_IWL<15595> A_IWL<15594> A_IWL<15593> A_IWL<15592> A_IWL<15591> A_IWL<15590> A_IWL<15589> A_IWL<15588> A_IWL<15587> A_IWL<15586> A_IWL<15585> A_IWL<15584> A_IWL<15583> A_IWL<15582> A_IWL<15581> A_IWL<15580> A_IWL<15579> A_IWL<15578> A_IWL<15577> A_IWL<15576> A_IWL<15575> A_IWL<15574> A_IWL<15573> A_IWL<15572> A_IWL<15571> A_IWL<15570> A_IWL<15569> A_IWL<15568> A_IWL<15567> A_IWL<15566> A_IWL<15565> A_IWL<15564> A_IWL<15563> A_IWL<15562> A_IWL<15561> A_IWL<15560> A_IWL<15559> A_IWL<15558> A_IWL<15557> A_IWL<15556> A_IWL<15555> A_IWL<15554> A_IWL<15553> A_IWL<15552> A_IWL<15551> A_IWL<15550> A_IWL<15549> A_IWL<15548> A_IWL<15547> A_IWL<15546> A_IWL<15545> A_IWL<15544> A_IWL<15543> A_IWL<15542> A_IWL<15541> A_IWL<15540> A_IWL<15539> A_IWL<15538> A_IWL<15537> A_IWL<15536> A_IWL<15535> A_IWL<15534> A_IWL<15533> A_IWL<15532> A_IWL<15531> A_IWL<15530> A_IWL<15529> A_IWL<15528> A_IWL<15527> A_IWL<15526> A_IWL<15525> A_IWL<15524> A_IWL<15523> A_IWL<15522> A_IWL<15521> A_IWL<15520> A_IWL<15519> A_IWL<15518> A_IWL<15517> A_IWL<15516> A_IWL<15515> A_IWL<15514> A_IWL<15513> A_IWL<15512> A_IWL<15511> A_IWL<15510> A_IWL<15509> A_IWL<15508> A_IWL<15507> A_IWL<15506> A_IWL<15505> A_IWL<15504> A_IWL<15503> A_IWL<15502> A_IWL<15501> A_IWL<15500> A_IWL<15499> A_IWL<15498> A_IWL<15497> A_IWL<15496> A_IWL<15495> A_IWL<15494> A_IWL<15493> A_IWL<15492> A_IWL<15491> A_IWL<15490> A_IWL<15489> A_IWL<15488> A_IWL<15487> A_IWL<15486> A_IWL<15485> A_IWL<15484> A_IWL<15483> A_IWL<15482> A_IWL<15481> A_IWL<15480> A_IWL<15479> A_IWL<15478> A_IWL<15477> A_IWL<15476> A_IWL<15475> A_IWL<15474> A_IWL<15473> A_IWL<15472> A_IWL<15471> A_IWL<15470> A_IWL<15469> A_IWL<15468> A_IWL<15467> A_IWL<15466> A_IWL<15465> A_IWL<15464> A_IWL<15463> A_IWL<15462> A_IWL<15461> A_IWL<15460> A_IWL<15459> A_IWL<15458> A_IWL<15457> A_IWL<15456> A_IWL<15455> A_IWL<15454> A_IWL<15453> A_IWL<15452> A_IWL<15451> A_IWL<15450> A_IWL<15449> A_IWL<15448> A_IWL<15447> A_IWL<15446> A_IWL<15445> A_IWL<15444> A_IWL<15443> A_IWL<15442> A_IWL<15441> A_IWL<15440> A_IWL<15439> A_IWL<15438> A_IWL<15437> A_IWL<15436> A_IWL<15435> A_IWL<15434> A_IWL<15433> A_IWL<15432> A_IWL<15431> A_IWL<15430> A_IWL<15429> A_IWL<15428> A_IWL<15427> A_IWL<15426> A_IWL<15425> A_IWL<15424> A_IWL<15423> A_IWL<15422> A_IWL<15421> A_IWL<15420> A_IWL<15419> A_IWL<15418> A_IWL<15417> A_IWL<15416> A_IWL<15415> A_IWL<15414> A_IWL<15413> A_IWL<15412> A_IWL<15411> A_IWL<15410> A_IWL<15409> A_IWL<15408> A_IWL<15407> A_IWL<15406> A_IWL<15405> A_IWL<15404> A_IWL<15403> A_IWL<15402> A_IWL<15401> A_IWL<15400> A_IWL<15399> A_IWL<15398> A_IWL<15397> A_IWL<15396> A_IWL<15395> A_IWL<15394> A_IWL<15393> A_IWL<15392> A_IWL<15391> A_IWL<15390> A_IWL<15389> A_IWL<15388> A_IWL<15387> A_IWL<15386> A_IWL<15385> A_IWL<15384> A_IWL<15383> A_IWL<15382> A_IWL<15381> A_IWL<15380> A_IWL<15379> A_IWL<15378> A_IWL<15377> A_IWL<15376> A_IWL<15375> A_IWL<15374> A_IWL<15373> A_IWL<15372> A_IWL<15371> A_IWL<15370> A_IWL<15369> A_IWL<15368> A_IWL<15367> A_IWL<15366> A_IWL<15365> A_IWL<15364> A_IWL<15363> A_IWL<15362> A_IWL<15361> A_IWL<15360> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<59> A_BLC<119> A_BLC<118> A_BLC_TOP<119> A_BLC_TOP<118> A_BLT<119> A_BLT<118> A_BLT_TOP<119> A_BLT_TOP<118> A_IWL<15103> A_IWL<15102> A_IWL<15101> A_IWL<15100> A_IWL<15099> A_IWL<15098> A_IWL<15097> A_IWL<15096> A_IWL<15095> A_IWL<15094> A_IWL<15093> A_IWL<15092> A_IWL<15091> A_IWL<15090> A_IWL<15089> A_IWL<15088> A_IWL<15087> A_IWL<15086> A_IWL<15085> A_IWL<15084> A_IWL<15083> A_IWL<15082> A_IWL<15081> A_IWL<15080> A_IWL<15079> A_IWL<15078> A_IWL<15077> A_IWL<15076> A_IWL<15075> A_IWL<15074> A_IWL<15073> A_IWL<15072> A_IWL<15071> A_IWL<15070> A_IWL<15069> A_IWL<15068> A_IWL<15067> A_IWL<15066> A_IWL<15065> A_IWL<15064> A_IWL<15063> A_IWL<15062> A_IWL<15061> A_IWL<15060> A_IWL<15059> A_IWL<15058> A_IWL<15057> A_IWL<15056> A_IWL<15055> A_IWL<15054> A_IWL<15053> A_IWL<15052> A_IWL<15051> A_IWL<15050> A_IWL<15049> A_IWL<15048> A_IWL<15047> A_IWL<15046> A_IWL<15045> A_IWL<15044> A_IWL<15043> A_IWL<15042> A_IWL<15041> A_IWL<15040> A_IWL<15039> A_IWL<15038> A_IWL<15037> A_IWL<15036> A_IWL<15035> A_IWL<15034> A_IWL<15033> A_IWL<15032> A_IWL<15031> A_IWL<15030> A_IWL<15029> A_IWL<15028> A_IWL<15027> A_IWL<15026> A_IWL<15025> A_IWL<15024> A_IWL<15023> A_IWL<15022> A_IWL<15021> A_IWL<15020> A_IWL<15019> A_IWL<15018> A_IWL<15017> A_IWL<15016> A_IWL<15015> A_IWL<15014> A_IWL<15013> A_IWL<15012> A_IWL<15011> A_IWL<15010> A_IWL<15009> A_IWL<15008> A_IWL<15007> A_IWL<15006> A_IWL<15005> A_IWL<15004> A_IWL<15003> A_IWL<15002> A_IWL<15001> A_IWL<15000> A_IWL<14999> A_IWL<14998> A_IWL<14997> A_IWL<14996> A_IWL<14995> A_IWL<14994> A_IWL<14993> A_IWL<14992> A_IWL<14991> A_IWL<14990> A_IWL<14989> A_IWL<14988> A_IWL<14987> A_IWL<14986> A_IWL<14985> A_IWL<14984> A_IWL<14983> A_IWL<14982> A_IWL<14981> A_IWL<14980> A_IWL<14979> A_IWL<14978> A_IWL<14977> A_IWL<14976> A_IWL<14975> A_IWL<14974> A_IWL<14973> A_IWL<14972> A_IWL<14971> A_IWL<14970> A_IWL<14969> A_IWL<14968> A_IWL<14967> A_IWL<14966> A_IWL<14965> A_IWL<14964> A_IWL<14963> A_IWL<14962> A_IWL<14961> A_IWL<14960> A_IWL<14959> A_IWL<14958> A_IWL<14957> A_IWL<14956> A_IWL<14955> A_IWL<14954> A_IWL<14953> A_IWL<14952> A_IWL<14951> A_IWL<14950> A_IWL<14949> A_IWL<14948> A_IWL<14947> A_IWL<14946> A_IWL<14945> A_IWL<14944> A_IWL<14943> A_IWL<14942> A_IWL<14941> A_IWL<14940> A_IWL<14939> A_IWL<14938> A_IWL<14937> A_IWL<14936> A_IWL<14935> A_IWL<14934> A_IWL<14933> A_IWL<14932> A_IWL<14931> A_IWL<14930> A_IWL<14929> A_IWL<14928> A_IWL<14927> A_IWL<14926> A_IWL<14925> A_IWL<14924> A_IWL<14923> A_IWL<14922> A_IWL<14921> A_IWL<14920> A_IWL<14919> A_IWL<14918> A_IWL<14917> A_IWL<14916> A_IWL<14915> A_IWL<14914> A_IWL<14913> A_IWL<14912> A_IWL<14911> A_IWL<14910> A_IWL<14909> A_IWL<14908> A_IWL<14907> A_IWL<14906> A_IWL<14905> A_IWL<14904> A_IWL<14903> A_IWL<14902> A_IWL<14901> A_IWL<14900> A_IWL<14899> A_IWL<14898> A_IWL<14897> A_IWL<14896> A_IWL<14895> A_IWL<14894> A_IWL<14893> A_IWL<14892> A_IWL<14891> A_IWL<14890> A_IWL<14889> A_IWL<14888> A_IWL<14887> A_IWL<14886> A_IWL<14885> A_IWL<14884> A_IWL<14883> A_IWL<14882> A_IWL<14881> A_IWL<14880> A_IWL<14879> A_IWL<14878> A_IWL<14877> A_IWL<14876> A_IWL<14875> A_IWL<14874> A_IWL<14873> A_IWL<14872> A_IWL<14871> A_IWL<14870> A_IWL<14869> A_IWL<14868> A_IWL<14867> A_IWL<14866> A_IWL<14865> A_IWL<14864> A_IWL<14863> A_IWL<14862> A_IWL<14861> A_IWL<14860> A_IWL<14859> A_IWL<14858> A_IWL<14857> A_IWL<14856> A_IWL<14855> A_IWL<14854> A_IWL<14853> A_IWL<14852> A_IWL<14851> A_IWL<14850> A_IWL<14849> A_IWL<14848> A_IWL<15359> A_IWL<15358> A_IWL<15357> A_IWL<15356> A_IWL<15355> A_IWL<15354> A_IWL<15353> A_IWL<15352> A_IWL<15351> A_IWL<15350> A_IWL<15349> A_IWL<15348> A_IWL<15347> A_IWL<15346> A_IWL<15345> A_IWL<15344> A_IWL<15343> A_IWL<15342> A_IWL<15341> A_IWL<15340> A_IWL<15339> A_IWL<15338> A_IWL<15337> A_IWL<15336> A_IWL<15335> A_IWL<15334> A_IWL<15333> A_IWL<15332> A_IWL<15331> A_IWL<15330> A_IWL<15329> A_IWL<15328> A_IWL<15327> A_IWL<15326> A_IWL<15325> A_IWL<15324> A_IWL<15323> A_IWL<15322> A_IWL<15321> A_IWL<15320> A_IWL<15319> A_IWL<15318> A_IWL<15317> A_IWL<15316> A_IWL<15315> A_IWL<15314> A_IWL<15313> A_IWL<15312> A_IWL<15311> A_IWL<15310> A_IWL<15309> A_IWL<15308> A_IWL<15307> A_IWL<15306> A_IWL<15305> A_IWL<15304> A_IWL<15303> A_IWL<15302> A_IWL<15301> A_IWL<15300> A_IWL<15299> A_IWL<15298> A_IWL<15297> A_IWL<15296> A_IWL<15295> A_IWL<15294> A_IWL<15293> A_IWL<15292> A_IWL<15291> A_IWL<15290> A_IWL<15289> A_IWL<15288> A_IWL<15287> A_IWL<15286> A_IWL<15285> A_IWL<15284> A_IWL<15283> A_IWL<15282> A_IWL<15281> A_IWL<15280> A_IWL<15279> A_IWL<15278> A_IWL<15277> A_IWL<15276> A_IWL<15275> A_IWL<15274> A_IWL<15273> A_IWL<15272> A_IWL<15271> A_IWL<15270> A_IWL<15269> A_IWL<15268> A_IWL<15267> A_IWL<15266> A_IWL<15265> A_IWL<15264> A_IWL<15263> A_IWL<15262> A_IWL<15261> A_IWL<15260> A_IWL<15259> A_IWL<15258> A_IWL<15257> A_IWL<15256> A_IWL<15255> A_IWL<15254> A_IWL<15253> A_IWL<15252> A_IWL<15251> A_IWL<15250> A_IWL<15249> A_IWL<15248> A_IWL<15247> A_IWL<15246> A_IWL<15245> A_IWL<15244> A_IWL<15243> A_IWL<15242> A_IWL<15241> A_IWL<15240> A_IWL<15239> A_IWL<15238> A_IWL<15237> A_IWL<15236> A_IWL<15235> A_IWL<15234> A_IWL<15233> A_IWL<15232> A_IWL<15231> A_IWL<15230> A_IWL<15229> A_IWL<15228> A_IWL<15227> A_IWL<15226> A_IWL<15225> A_IWL<15224> A_IWL<15223> A_IWL<15222> A_IWL<15221> A_IWL<15220> A_IWL<15219> A_IWL<15218> A_IWL<15217> A_IWL<15216> A_IWL<15215> A_IWL<15214> A_IWL<15213> A_IWL<15212> A_IWL<15211> A_IWL<15210> A_IWL<15209> A_IWL<15208> A_IWL<15207> A_IWL<15206> A_IWL<15205> A_IWL<15204> A_IWL<15203> A_IWL<15202> A_IWL<15201> A_IWL<15200> A_IWL<15199> A_IWL<15198> A_IWL<15197> A_IWL<15196> A_IWL<15195> A_IWL<15194> A_IWL<15193> A_IWL<15192> A_IWL<15191> A_IWL<15190> A_IWL<15189> A_IWL<15188> A_IWL<15187> A_IWL<15186> A_IWL<15185> A_IWL<15184> A_IWL<15183> A_IWL<15182> A_IWL<15181> A_IWL<15180> A_IWL<15179> A_IWL<15178> A_IWL<15177> A_IWL<15176> A_IWL<15175> A_IWL<15174> A_IWL<15173> A_IWL<15172> A_IWL<15171> A_IWL<15170> A_IWL<15169> A_IWL<15168> A_IWL<15167> A_IWL<15166> A_IWL<15165> A_IWL<15164> A_IWL<15163> A_IWL<15162> A_IWL<15161> A_IWL<15160> A_IWL<15159> A_IWL<15158> A_IWL<15157> A_IWL<15156> A_IWL<15155> A_IWL<15154> A_IWL<15153> A_IWL<15152> A_IWL<15151> A_IWL<15150> A_IWL<15149> A_IWL<15148> A_IWL<15147> A_IWL<15146> A_IWL<15145> A_IWL<15144> A_IWL<15143> A_IWL<15142> A_IWL<15141> A_IWL<15140> A_IWL<15139> A_IWL<15138> A_IWL<15137> A_IWL<15136> A_IWL<15135> A_IWL<15134> A_IWL<15133> A_IWL<15132> A_IWL<15131> A_IWL<15130> A_IWL<15129> A_IWL<15128> A_IWL<15127> A_IWL<15126> A_IWL<15125> A_IWL<15124> A_IWL<15123> A_IWL<15122> A_IWL<15121> A_IWL<15120> A_IWL<15119> A_IWL<15118> A_IWL<15117> A_IWL<15116> A_IWL<15115> A_IWL<15114> A_IWL<15113> A_IWL<15112> A_IWL<15111> A_IWL<15110> A_IWL<15109> A_IWL<15108> A_IWL<15107> A_IWL<15106> A_IWL<15105> A_IWL<15104> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<58> A_BLC<117> A_BLC<116> A_BLC_TOP<117> A_BLC_TOP<116> A_BLT<117> A_BLT<116> A_BLT_TOP<117> A_BLT_TOP<116> A_IWL<14847> A_IWL<14846> A_IWL<14845> A_IWL<14844> A_IWL<14843> A_IWL<14842> A_IWL<14841> A_IWL<14840> A_IWL<14839> A_IWL<14838> A_IWL<14837> A_IWL<14836> A_IWL<14835> A_IWL<14834> A_IWL<14833> A_IWL<14832> A_IWL<14831> A_IWL<14830> A_IWL<14829> A_IWL<14828> A_IWL<14827> A_IWL<14826> A_IWL<14825> A_IWL<14824> A_IWL<14823> A_IWL<14822> A_IWL<14821> A_IWL<14820> A_IWL<14819> A_IWL<14818> A_IWL<14817> A_IWL<14816> A_IWL<14815> A_IWL<14814> A_IWL<14813> A_IWL<14812> A_IWL<14811> A_IWL<14810> A_IWL<14809> A_IWL<14808> A_IWL<14807> A_IWL<14806> A_IWL<14805> A_IWL<14804> A_IWL<14803> A_IWL<14802> A_IWL<14801> A_IWL<14800> A_IWL<14799> A_IWL<14798> A_IWL<14797> A_IWL<14796> A_IWL<14795> A_IWL<14794> A_IWL<14793> A_IWL<14792> A_IWL<14791> A_IWL<14790> A_IWL<14789> A_IWL<14788> A_IWL<14787> A_IWL<14786> A_IWL<14785> A_IWL<14784> A_IWL<14783> A_IWL<14782> A_IWL<14781> A_IWL<14780> A_IWL<14779> A_IWL<14778> A_IWL<14777> A_IWL<14776> A_IWL<14775> A_IWL<14774> A_IWL<14773> A_IWL<14772> A_IWL<14771> A_IWL<14770> A_IWL<14769> A_IWL<14768> A_IWL<14767> A_IWL<14766> A_IWL<14765> A_IWL<14764> A_IWL<14763> A_IWL<14762> A_IWL<14761> A_IWL<14760> A_IWL<14759> A_IWL<14758> A_IWL<14757> A_IWL<14756> A_IWL<14755> A_IWL<14754> A_IWL<14753> A_IWL<14752> A_IWL<14751> A_IWL<14750> A_IWL<14749> A_IWL<14748> A_IWL<14747> A_IWL<14746> A_IWL<14745> A_IWL<14744> A_IWL<14743> A_IWL<14742> A_IWL<14741> A_IWL<14740> A_IWL<14739> A_IWL<14738> A_IWL<14737> A_IWL<14736> A_IWL<14735> A_IWL<14734> A_IWL<14733> A_IWL<14732> A_IWL<14731> A_IWL<14730> A_IWL<14729> A_IWL<14728> A_IWL<14727> A_IWL<14726> A_IWL<14725> A_IWL<14724> A_IWL<14723> A_IWL<14722> A_IWL<14721> A_IWL<14720> A_IWL<14719> A_IWL<14718> A_IWL<14717> A_IWL<14716> A_IWL<14715> A_IWL<14714> A_IWL<14713> A_IWL<14712> A_IWL<14711> A_IWL<14710> A_IWL<14709> A_IWL<14708> A_IWL<14707> A_IWL<14706> A_IWL<14705> A_IWL<14704> A_IWL<14703> A_IWL<14702> A_IWL<14701> A_IWL<14700> A_IWL<14699> A_IWL<14698> A_IWL<14697> A_IWL<14696> A_IWL<14695> A_IWL<14694> A_IWL<14693> A_IWL<14692> A_IWL<14691> A_IWL<14690> A_IWL<14689> A_IWL<14688> A_IWL<14687> A_IWL<14686> A_IWL<14685> A_IWL<14684> A_IWL<14683> A_IWL<14682> A_IWL<14681> A_IWL<14680> A_IWL<14679> A_IWL<14678> A_IWL<14677> A_IWL<14676> A_IWL<14675> A_IWL<14674> A_IWL<14673> A_IWL<14672> A_IWL<14671> A_IWL<14670> A_IWL<14669> A_IWL<14668> A_IWL<14667> A_IWL<14666> A_IWL<14665> A_IWL<14664> A_IWL<14663> A_IWL<14662> A_IWL<14661> A_IWL<14660> A_IWL<14659> A_IWL<14658> A_IWL<14657> A_IWL<14656> A_IWL<14655> A_IWL<14654> A_IWL<14653> A_IWL<14652> A_IWL<14651> A_IWL<14650> A_IWL<14649> A_IWL<14648> A_IWL<14647> A_IWL<14646> A_IWL<14645> A_IWL<14644> A_IWL<14643> A_IWL<14642> A_IWL<14641> A_IWL<14640> A_IWL<14639> A_IWL<14638> A_IWL<14637> A_IWL<14636> A_IWL<14635> A_IWL<14634> A_IWL<14633> A_IWL<14632> A_IWL<14631> A_IWL<14630> A_IWL<14629> A_IWL<14628> A_IWL<14627> A_IWL<14626> A_IWL<14625> A_IWL<14624> A_IWL<14623> A_IWL<14622> A_IWL<14621> A_IWL<14620> A_IWL<14619> A_IWL<14618> A_IWL<14617> A_IWL<14616> A_IWL<14615> A_IWL<14614> A_IWL<14613> A_IWL<14612> A_IWL<14611> A_IWL<14610> A_IWL<14609> A_IWL<14608> A_IWL<14607> A_IWL<14606> A_IWL<14605> A_IWL<14604> A_IWL<14603> A_IWL<14602> A_IWL<14601> A_IWL<14600> A_IWL<14599> A_IWL<14598> A_IWL<14597> A_IWL<14596> A_IWL<14595> A_IWL<14594> A_IWL<14593> A_IWL<14592> A_IWL<15103> A_IWL<15102> A_IWL<15101> A_IWL<15100> A_IWL<15099> A_IWL<15098> A_IWL<15097> A_IWL<15096> A_IWL<15095> A_IWL<15094> A_IWL<15093> A_IWL<15092> A_IWL<15091> A_IWL<15090> A_IWL<15089> A_IWL<15088> A_IWL<15087> A_IWL<15086> A_IWL<15085> A_IWL<15084> A_IWL<15083> A_IWL<15082> A_IWL<15081> A_IWL<15080> A_IWL<15079> A_IWL<15078> A_IWL<15077> A_IWL<15076> A_IWL<15075> A_IWL<15074> A_IWL<15073> A_IWL<15072> A_IWL<15071> A_IWL<15070> A_IWL<15069> A_IWL<15068> A_IWL<15067> A_IWL<15066> A_IWL<15065> A_IWL<15064> A_IWL<15063> A_IWL<15062> A_IWL<15061> A_IWL<15060> A_IWL<15059> A_IWL<15058> A_IWL<15057> A_IWL<15056> A_IWL<15055> A_IWL<15054> A_IWL<15053> A_IWL<15052> A_IWL<15051> A_IWL<15050> A_IWL<15049> A_IWL<15048> A_IWL<15047> A_IWL<15046> A_IWL<15045> A_IWL<15044> A_IWL<15043> A_IWL<15042> A_IWL<15041> A_IWL<15040> A_IWL<15039> A_IWL<15038> A_IWL<15037> A_IWL<15036> A_IWL<15035> A_IWL<15034> A_IWL<15033> A_IWL<15032> A_IWL<15031> A_IWL<15030> A_IWL<15029> A_IWL<15028> A_IWL<15027> A_IWL<15026> A_IWL<15025> A_IWL<15024> A_IWL<15023> A_IWL<15022> A_IWL<15021> A_IWL<15020> A_IWL<15019> A_IWL<15018> A_IWL<15017> A_IWL<15016> A_IWL<15015> A_IWL<15014> A_IWL<15013> A_IWL<15012> A_IWL<15011> A_IWL<15010> A_IWL<15009> A_IWL<15008> A_IWL<15007> A_IWL<15006> A_IWL<15005> A_IWL<15004> A_IWL<15003> A_IWL<15002> A_IWL<15001> A_IWL<15000> A_IWL<14999> A_IWL<14998> A_IWL<14997> A_IWL<14996> A_IWL<14995> A_IWL<14994> A_IWL<14993> A_IWL<14992> A_IWL<14991> A_IWL<14990> A_IWL<14989> A_IWL<14988> A_IWL<14987> A_IWL<14986> A_IWL<14985> A_IWL<14984> A_IWL<14983> A_IWL<14982> A_IWL<14981> A_IWL<14980> A_IWL<14979> A_IWL<14978> A_IWL<14977> A_IWL<14976> A_IWL<14975> A_IWL<14974> A_IWL<14973> A_IWL<14972> A_IWL<14971> A_IWL<14970> A_IWL<14969> A_IWL<14968> A_IWL<14967> A_IWL<14966> A_IWL<14965> A_IWL<14964> A_IWL<14963> A_IWL<14962> A_IWL<14961> A_IWL<14960> A_IWL<14959> A_IWL<14958> A_IWL<14957> A_IWL<14956> A_IWL<14955> A_IWL<14954> A_IWL<14953> A_IWL<14952> A_IWL<14951> A_IWL<14950> A_IWL<14949> A_IWL<14948> A_IWL<14947> A_IWL<14946> A_IWL<14945> A_IWL<14944> A_IWL<14943> A_IWL<14942> A_IWL<14941> A_IWL<14940> A_IWL<14939> A_IWL<14938> A_IWL<14937> A_IWL<14936> A_IWL<14935> A_IWL<14934> A_IWL<14933> A_IWL<14932> A_IWL<14931> A_IWL<14930> A_IWL<14929> A_IWL<14928> A_IWL<14927> A_IWL<14926> A_IWL<14925> A_IWL<14924> A_IWL<14923> A_IWL<14922> A_IWL<14921> A_IWL<14920> A_IWL<14919> A_IWL<14918> A_IWL<14917> A_IWL<14916> A_IWL<14915> A_IWL<14914> A_IWL<14913> A_IWL<14912> A_IWL<14911> A_IWL<14910> A_IWL<14909> A_IWL<14908> A_IWL<14907> A_IWL<14906> A_IWL<14905> A_IWL<14904> A_IWL<14903> A_IWL<14902> A_IWL<14901> A_IWL<14900> A_IWL<14899> A_IWL<14898> A_IWL<14897> A_IWL<14896> A_IWL<14895> A_IWL<14894> A_IWL<14893> A_IWL<14892> A_IWL<14891> A_IWL<14890> A_IWL<14889> A_IWL<14888> A_IWL<14887> A_IWL<14886> A_IWL<14885> A_IWL<14884> A_IWL<14883> A_IWL<14882> A_IWL<14881> A_IWL<14880> A_IWL<14879> A_IWL<14878> A_IWL<14877> A_IWL<14876> A_IWL<14875> A_IWL<14874> A_IWL<14873> A_IWL<14872> A_IWL<14871> A_IWL<14870> A_IWL<14869> A_IWL<14868> A_IWL<14867> A_IWL<14866> A_IWL<14865> A_IWL<14864> A_IWL<14863> A_IWL<14862> A_IWL<14861> A_IWL<14860> A_IWL<14859> A_IWL<14858> A_IWL<14857> A_IWL<14856> A_IWL<14855> A_IWL<14854> A_IWL<14853> A_IWL<14852> A_IWL<14851> A_IWL<14850> A_IWL<14849> A_IWL<14848> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<57> A_BLC<115> A_BLC<114> A_BLC_TOP<115> A_BLC_TOP<114> A_BLT<115> A_BLT<114> A_BLT_TOP<115> A_BLT_TOP<114> A_IWL<14591> A_IWL<14590> A_IWL<14589> A_IWL<14588> A_IWL<14587> A_IWL<14586> A_IWL<14585> A_IWL<14584> A_IWL<14583> A_IWL<14582> A_IWL<14581> A_IWL<14580> A_IWL<14579> A_IWL<14578> A_IWL<14577> A_IWL<14576> A_IWL<14575> A_IWL<14574> A_IWL<14573> A_IWL<14572> A_IWL<14571> A_IWL<14570> A_IWL<14569> A_IWL<14568> A_IWL<14567> A_IWL<14566> A_IWL<14565> A_IWL<14564> A_IWL<14563> A_IWL<14562> A_IWL<14561> A_IWL<14560> A_IWL<14559> A_IWL<14558> A_IWL<14557> A_IWL<14556> A_IWL<14555> A_IWL<14554> A_IWL<14553> A_IWL<14552> A_IWL<14551> A_IWL<14550> A_IWL<14549> A_IWL<14548> A_IWL<14547> A_IWL<14546> A_IWL<14545> A_IWL<14544> A_IWL<14543> A_IWL<14542> A_IWL<14541> A_IWL<14540> A_IWL<14539> A_IWL<14538> A_IWL<14537> A_IWL<14536> A_IWL<14535> A_IWL<14534> A_IWL<14533> A_IWL<14532> A_IWL<14531> A_IWL<14530> A_IWL<14529> A_IWL<14528> A_IWL<14527> A_IWL<14526> A_IWL<14525> A_IWL<14524> A_IWL<14523> A_IWL<14522> A_IWL<14521> A_IWL<14520> A_IWL<14519> A_IWL<14518> A_IWL<14517> A_IWL<14516> A_IWL<14515> A_IWL<14514> A_IWL<14513> A_IWL<14512> A_IWL<14511> A_IWL<14510> A_IWL<14509> A_IWL<14508> A_IWL<14507> A_IWL<14506> A_IWL<14505> A_IWL<14504> A_IWL<14503> A_IWL<14502> A_IWL<14501> A_IWL<14500> A_IWL<14499> A_IWL<14498> A_IWL<14497> A_IWL<14496> A_IWL<14495> A_IWL<14494> A_IWL<14493> A_IWL<14492> A_IWL<14491> A_IWL<14490> A_IWL<14489> A_IWL<14488> A_IWL<14487> A_IWL<14486> A_IWL<14485> A_IWL<14484> A_IWL<14483> A_IWL<14482> A_IWL<14481> A_IWL<14480> A_IWL<14479> A_IWL<14478> A_IWL<14477> A_IWL<14476> A_IWL<14475> A_IWL<14474> A_IWL<14473> A_IWL<14472> A_IWL<14471> A_IWL<14470> A_IWL<14469> A_IWL<14468> A_IWL<14467> A_IWL<14466> A_IWL<14465> A_IWL<14464> A_IWL<14463> A_IWL<14462> A_IWL<14461> A_IWL<14460> A_IWL<14459> A_IWL<14458> A_IWL<14457> A_IWL<14456> A_IWL<14455> A_IWL<14454> A_IWL<14453> A_IWL<14452> A_IWL<14451> A_IWL<14450> A_IWL<14449> A_IWL<14448> A_IWL<14447> A_IWL<14446> A_IWL<14445> A_IWL<14444> A_IWL<14443> A_IWL<14442> A_IWL<14441> A_IWL<14440> A_IWL<14439> A_IWL<14438> A_IWL<14437> A_IWL<14436> A_IWL<14435> A_IWL<14434> A_IWL<14433> A_IWL<14432> A_IWL<14431> A_IWL<14430> A_IWL<14429> A_IWL<14428> A_IWL<14427> A_IWL<14426> A_IWL<14425> A_IWL<14424> A_IWL<14423> A_IWL<14422> A_IWL<14421> A_IWL<14420> A_IWL<14419> A_IWL<14418> A_IWL<14417> A_IWL<14416> A_IWL<14415> A_IWL<14414> A_IWL<14413> A_IWL<14412> A_IWL<14411> A_IWL<14410> A_IWL<14409> A_IWL<14408> A_IWL<14407> A_IWL<14406> A_IWL<14405> A_IWL<14404> A_IWL<14403> A_IWL<14402> A_IWL<14401> A_IWL<14400> A_IWL<14399> A_IWL<14398> A_IWL<14397> A_IWL<14396> A_IWL<14395> A_IWL<14394> A_IWL<14393> A_IWL<14392> A_IWL<14391> A_IWL<14390> A_IWL<14389> A_IWL<14388> A_IWL<14387> A_IWL<14386> A_IWL<14385> A_IWL<14384> A_IWL<14383> A_IWL<14382> A_IWL<14381> A_IWL<14380> A_IWL<14379> A_IWL<14378> A_IWL<14377> A_IWL<14376> A_IWL<14375> A_IWL<14374> A_IWL<14373> A_IWL<14372> A_IWL<14371> A_IWL<14370> A_IWL<14369> A_IWL<14368> A_IWL<14367> A_IWL<14366> A_IWL<14365> A_IWL<14364> A_IWL<14363> A_IWL<14362> A_IWL<14361> A_IWL<14360> A_IWL<14359> A_IWL<14358> A_IWL<14357> A_IWL<14356> A_IWL<14355> A_IWL<14354> A_IWL<14353> A_IWL<14352> A_IWL<14351> A_IWL<14350> A_IWL<14349> A_IWL<14348> A_IWL<14347> A_IWL<14346> A_IWL<14345> A_IWL<14344> A_IWL<14343> A_IWL<14342> A_IWL<14341> A_IWL<14340> A_IWL<14339> A_IWL<14338> A_IWL<14337> A_IWL<14336> A_IWL<14847> A_IWL<14846> A_IWL<14845> A_IWL<14844> A_IWL<14843> A_IWL<14842> A_IWL<14841> A_IWL<14840> A_IWL<14839> A_IWL<14838> A_IWL<14837> A_IWL<14836> A_IWL<14835> A_IWL<14834> A_IWL<14833> A_IWL<14832> A_IWL<14831> A_IWL<14830> A_IWL<14829> A_IWL<14828> A_IWL<14827> A_IWL<14826> A_IWL<14825> A_IWL<14824> A_IWL<14823> A_IWL<14822> A_IWL<14821> A_IWL<14820> A_IWL<14819> A_IWL<14818> A_IWL<14817> A_IWL<14816> A_IWL<14815> A_IWL<14814> A_IWL<14813> A_IWL<14812> A_IWL<14811> A_IWL<14810> A_IWL<14809> A_IWL<14808> A_IWL<14807> A_IWL<14806> A_IWL<14805> A_IWL<14804> A_IWL<14803> A_IWL<14802> A_IWL<14801> A_IWL<14800> A_IWL<14799> A_IWL<14798> A_IWL<14797> A_IWL<14796> A_IWL<14795> A_IWL<14794> A_IWL<14793> A_IWL<14792> A_IWL<14791> A_IWL<14790> A_IWL<14789> A_IWL<14788> A_IWL<14787> A_IWL<14786> A_IWL<14785> A_IWL<14784> A_IWL<14783> A_IWL<14782> A_IWL<14781> A_IWL<14780> A_IWL<14779> A_IWL<14778> A_IWL<14777> A_IWL<14776> A_IWL<14775> A_IWL<14774> A_IWL<14773> A_IWL<14772> A_IWL<14771> A_IWL<14770> A_IWL<14769> A_IWL<14768> A_IWL<14767> A_IWL<14766> A_IWL<14765> A_IWL<14764> A_IWL<14763> A_IWL<14762> A_IWL<14761> A_IWL<14760> A_IWL<14759> A_IWL<14758> A_IWL<14757> A_IWL<14756> A_IWL<14755> A_IWL<14754> A_IWL<14753> A_IWL<14752> A_IWL<14751> A_IWL<14750> A_IWL<14749> A_IWL<14748> A_IWL<14747> A_IWL<14746> A_IWL<14745> A_IWL<14744> A_IWL<14743> A_IWL<14742> A_IWL<14741> A_IWL<14740> A_IWL<14739> A_IWL<14738> A_IWL<14737> A_IWL<14736> A_IWL<14735> A_IWL<14734> A_IWL<14733> A_IWL<14732> A_IWL<14731> A_IWL<14730> A_IWL<14729> A_IWL<14728> A_IWL<14727> A_IWL<14726> A_IWL<14725> A_IWL<14724> A_IWL<14723> A_IWL<14722> A_IWL<14721> A_IWL<14720> A_IWL<14719> A_IWL<14718> A_IWL<14717> A_IWL<14716> A_IWL<14715> A_IWL<14714> A_IWL<14713> A_IWL<14712> A_IWL<14711> A_IWL<14710> A_IWL<14709> A_IWL<14708> A_IWL<14707> A_IWL<14706> A_IWL<14705> A_IWL<14704> A_IWL<14703> A_IWL<14702> A_IWL<14701> A_IWL<14700> A_IWL<14699> A_IWL<14698> A_IWL<14697> A_IWL<14696> A_IWL<14695> A_IWL<14694> A_IWL<14693> A_IWL<14692> A_IWL<14691> A_IWL<14690> A_IWL<14689> A_IWL<14688> A_IWL<14687> A_IWL<14686> A_IWL<14685> A_IWL<14684> A_IWL<14683> A_IWL<14682> A_IWL<14681> A_IWL<14680> A_IWL<14679> A_IWL<14678> A_IWL<14677> A_IWL<14676> A_IWL<14675> A_IWL<14674> A_IWL<14673> A_IWL<14672> A_IWL<14671> A_IWL<14670> A_IWL<14669> A_IWL<14668> A_IWL<14667> A_IWL<14666> A_IWL<14665> A_IWL<14664> A_IWL<14663> A_IWL<14662> A_IWL<14661> A_IWL<14660> A_IWL<14659> A_IWL<14658> A_IWL<14657> A_IWL<14656> A_IWL<14655> A_IWL<14654> A_IWL<14653> A_IWL<14652> A_IWL<14651> A_IWL<14650> A_IWL<14649> A_IWL<14648> A_IWL<14647> A_IWL<14646> A_IWL<14645> A_IWL<14644> A_IWL<14643> A_IWL<14642> A_IWL<14641> A_IWL<14640> A_IWL<14639> A_IWL<14638> A_IWL<14637> A_IWL<14636> A_IWL<14635> A_IWL<14634> A_IWL<14633> A_IWL<14632> A_IWL<14631> A_IWL<14630> A_IWL<14629> A_IWL<14628> A_IWL<14627> A_IWL<14626> A_IWL<14625> A_IWL<14624> A_IWL<14623> A_IWL<14622> A_IWL<14621> A_IWL<14620> A_IWL<14619> A_IWL<14618> A_IWL<14617> A_IWL<14616> A_IWL<14615> A_IWL<14614> A_IWL<14613> A_IWL<14612> A_IWL<14611> A_IWL<14610> A_IWL<14609> A_IWL<14608> A_IWL<14607> A_IWL<14606> A_IWL<14605> A_IWL<14604> A_IWL<14603> A_IWL<14602> A_IWL<14601> A_IWL<14600> A_IWL<14599> A_IWL<14598> A_IWL<14597> A_IWL<14596> A_IWL<14595> A_IWL<14594> A_IWL<14593> A_IWL<14592> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<56> A_BLC<113> A_BLC<112> A_BLC_TOP<113> A_BLC_TOP<112> A_BLT<113> A_BLT<112> A_BLT_TOP<113> A_BLT_TOP<112> A_IWL<14335> A_IWL<14334> A_IWL<14333> A_IWL<14332> A_IWL<14331> A_IWL<14330> A_IWL<14329> A_IWL<14328> A_IWL<14327> A_IWL<14326> A_IWL<14325> A_IWL<14324> A_IWL<14323> A_IWL<14322> A_IWL<14321> A_IWL<14320> A_IWL<14319> A_IWL<14318> A_IWL<14317> A_IWL<14316> A_IWL<14315> A_IWL<14314> A_IWL<14313> A_IWL<14312> A_IWL<14311> A_IWL<14310> A_IWL<14309> A_IWL<14308> A_IWL<14307> A_IWL<14306> A_IWL<14305> A_IWL<14304> A_IWL<14303> A_IWL<14302> A_IWL<14301> A_IWL<14300> A_IWL<14299> A_IWL<14298> A_IWL<14297> A_IWL<14296> A_IWL<14295> A_IWL<14294> A_IWL<14293> A_IWL<14292> A_IWL<14291> A_IWL<14290> A_IWL<14289> A_IWL<14288> A_IWL<14287> A_IWL<14286> A_IWL<14285> A_IWL<14284> A_IWL<14283> A_IWL<14282> A_IWL<14281> A_IWL<14280> A_IWL<14279> A_IWL<14278> A_IWL<14277> A_IWL<14276> A_IWL<14275> A_IWL<14274> A_IWL<14273> A_IWL<14272> A_IWL<14271> A_IWL<14270> A_IWL<14269> A_IWL<14268> A_IWL<14267> A_IWL<14266> A_IWL<14265> A_IWL<14264> A_IWL<14263> A_IWL<14262> A_IWL<14261> A_IWL<14260> A_IWL<14259> A_IWL<14258> A_IWL<14257> A_IWL<14256> A_IWL<14255> A_IWL<14254> A_IWL<14253> A_IWL<14252> A_IWL<14251> A_IWL<14250> A_IWL<14249> A_IWL<14248> A_IWL<14247> A_IWL<14246> A_IWL<14245> A_IWL<14244> A_IWL<14243> A_IWL<14242> A_IWL<14241> A_IWL<14240> A_IWL<14239> A_IWL<14238> A_IWL<14237> A_IWL<14236> A_IWL<14235> A_IWL<14234> A_IWL<14233> A_IWL<14232> A_IWL<14231> A_IWL<14230> A_IWL<14229> A_IWL<14228> A_IWL<14227> A_IWL<14226> A_IWL<14225> A_IWL<14224> A_IWL<14223> A_IWL<14222> A_IWL<14221> A_IWL<14220> A_IWL<14219> A_IWL<14218> A_IWL<14217> A_IWL<14216> A_IWL<14215> A_IWL<14214> A_IWL<14213> A_IWL<14212> A_IWL<14211> A_IWL<14210> A_IWL<14209> A_IWL<14208> A_IWL<14207> A_IWL<14206> A_IWL<14205> A_IWL<14204> A_IWL<14203> A_IWL<14202> A_IWL<14201> A_IWL<14200> A_IWL<14199> A_IWL<14198> A_IWL<14197> A_IWL<14196> A_IWL<14195> A_IWL<14194> A_IWL<14193> A_IWL<14192> A_IWL<14191> A_IWL<14190> A_IWL<14189> A_IWL<14188> A_IWL<14187> A_IWL<14186> A_IWL<14185> A_IWL<14184> A_IWL<14183> A_IWL<14182> A_IWL<14181> A_IWL<14180> A_IWL<14179> A_IWL<14178> A_IWL<14177> A_IWL<14176> A_IWL<14175> A_IWL<14174> A_IWL<14173> A_IWL<14172> A_IWL<14171> A_IWL<14170> A_IWL<14169> A_IWL<14168> A_IWL<14167> A_IWL<14166> A_IWL<14165> A_IWL<14164> A_IWL<14163> A_IWL<14162> A_IWL<14161> A_IWL<14160> A_IWL<14159> A_IWL<14158> A_IWL<14157> A_IWL<14156> A_IWL<14155> A_IWL<14154> A_IWL<14153> A_IWL<14152> A_IWL<14151> A_IWL<14150> A_IWL<14149> A_IWL<14148> A_IWL<14147> A_IWL<14146> A_IWL<14145> A_IWL<14144> A_IWL<14143> A_IWL<14142> A_IWL<14141> A_IWL<14140> A_IWL<14139> A_IWL<14138> A_IWL<14137> A_IWL<14136> A_IWL<14135> A_IWL<14134> A_IWL<14133> A_IWL<14132> A_IWL<14131> A_IWL<14130> A_IWL<14129> A_IWL<14128> A_IWL<14127> A_IWL<14126> A_IWL<14125> A_IWL<14124> A_IWL<14123> A_IWL<14122> A_IWL<14121> A_IWL<14120> A_IWL<14119> A_IWL<14118> A_IWL<14117> A_IWL<14116> A_IWL<14115> A_IWL<14114> A_IWL<14113> A_IWL<14112> A_IWL<14111> A_IWL<14110> A_IWL<14109> A_IWL<14108> A_IWL<14107> A_IWL<14106> A_IWL<14105> A_IWL<14104> A_IWL<14103> A_IWL<14102> A_IWL<14101> A_IWL<14100> A_IWL<14099> A_IWL<14098> A_IWL<14097> A_IWL<14096> A_IWL<14095> A_IWL<14094> A_IWL<14093> A_IWL<14092> A_IWL<14091> A_IWL<14090> A_IWL<14089> A_IWL<14088> A_IWL<14087> A_IWL<14086> A_IWL<14085> A_IWL<14084> A_IWL<14083> A_IWL<14082> A_IWL<14081> A_IWL<14080> A_IWL<14591> A_IWL<14590> A_IWL<14589> A_IWL<14588> A_IWL<14587> A_IWL<14586> A_IWL<14585> A_IWL<14584> A_IWL<14583> A_IWL<14582> A_IWL<14581> A_IWL<14580> A_IWL<14579> A_IWL<14578> A_IWL<14577> A_IWL<14576> A_IWL<14575> A_IWL<14574> A_IWL<14573> A_IWL<14572> A_IWL<14571> A_IWL<14570> A_IWL<14569> A_IWL<14568> A_IWL<14567> A_IWL<14566> A_IWL<14565> A_IWL<14564> A_IWL<14563> A_IWL<14562> A_IWL<14561> A_IWL<14560> A_IWL<14559> A_IWL<14558> A_IWL<14557> A_IWL<14556> A_IWL<14555> A_IWL<14554> A_IWL<14553> A_IWL<14552> A_IWL<14551> A_IWL<14550> A_IWL<14549> A_IWL<14548> A_IWL<14547> A_IWL<14546> A_IWL<14545> A_IWL<14544> A_IWL<14543> A_IWL<14542> A_IWL<14541> A_IWL<14540> A_IWL<14539> A_IWL<14538> A_IWL<14537> A_IWL<14536> A_IWL<14535> A_IWL<14534> A_IWL<14533> A_IWL<14532> A_IWL<14531> A_IWL<14530> A_IWL<14529> A_IWL<14528> A_IWL<14527> A_IWL<14526> A_IWL<14525> A_IWL<14524> A_IWL<14523> A_IWL<14522> A_IWL<14521> A_IWL<14520> A_IWL<14519> A_IWL<14518> A_IWL<14517> A_IWL<14516> A_IWL<14515> A_IWL<14514> A_IWL<14513> A_IWL<14512> A_IWL<14511> A_IWL<14510> A_IWL<14509> A_IWL<14508> A_IWL<14507> A_IWL<14506> A_IWL<14505> A_IWL<14504> A_IWL<14503> A_IWL<14502> A_IWL<14501> A_IWL<14500> A_IWL<14499> A_IWL<14498> A_IWL<14497> A_IWL<14496> A_IWL<14495> A_IWL<14494> A_IWL<14493> A_IWL<14492> A_IWL<14491> A_IWL<14490> A_IWL<14489> A_IWL<14488> A_IWL<14487> A_IWL<14486> A_IWL<14485> A_IWL<14484> A_IWL<14483> A_IWL<14482> A_IWL<14481> A_IWL<14480> A_IWL<14479> A_IWL<14478> A_IWL<14477> A_IWL<14476> A_IWL<14475> A_IWL<14474> A_IWL<14473> A_IWL<14472> A_IWL<14471> A_IWL<14470> A_IWL<14469> A_IWL<14468> A_IWL<14467> A_IWL<14466> A_IWL<14465> A_IWL<14464> A_IWL<14463> A_IWL<14462> A_IWL<14461> A_IWL<14460> A_IWL<14459> A_IWL<14458> A_IWL<14457> A_IWL<14456> A_IWL<14455> A_IWL<14454> A_IWL<14453> A_IWL<14452> A_IWL<14451> A_IWL<14450> A_IWL<14449> A_IWL<14448> A_IWL<14447> A_IWL<14446> A_IWL<14445> A_IWL<14444> A_IWL<14443> A_IWL<14442> A_IWL<14441> A_IWL<14440> A_IWL<14439> A_IWL<14438> A_IWL<14437> A_IWL<14436> A_IWL<14435> A_IWL<14434> A_IWL<14433> A_IWL<14432> A_IWL<14431> A_IWL<14430> A_IWL<14429> A_IWL<14428> A_IWL<14427> A_IWL<14426> A_IWL<14425> A_IWL<14424> A_IWL<14423> A_IWL<14422> A_IWL<14421> A_IWL<14420> A_IWL<14419> A_IWL<14418> A_IWL<14417> A_IWL<14416> A_IWL<14415> A_IWL<14414> A_IWL<14413> A_IWL<14412> A_IWL<14411> A_IWL<14410> A_IWL<14409> A_IWL<14408> A_IWL<14407> A_IWL<14406> A_IWL<14405> A_IWL<14404> A_IWL<14403> A_IWL<14402> A_IWL<14401> A_IWL<14400> A_IWL<14399> A_IWL<14398> A_IWL<14397> A_IWL<14396> A_IWL<14395> A_IWL<14394> A_IWL<14393> A_IWL<14392> A_IWL<14391> A_IWL<14390> A_IWL<14389> A_IWL<14388> A_IWL<14387> A_IWL<14386> A_IWL<14385> A_IWL<14384> A_IWL<14383> A_IWL<14382> A_IWL<14381> A_IWL<14380> A_IWL<14379> A_IWL<14378> A_IWL<14377> A_IWL<14376> A_IWL<14375> A_IWL<14374> A_IWL<14373> A_IWL<14372> A_IWL<14371> A_IWL<14370> A_IWL<14369> A_IWL<14368> A_IWL<14367> A_IWL<14366> A_IWL<14365> A_IWL<14364> A_IWL<14363> A_IWL<14362> A_IWL<14361> A_IWL<14360> A_IWL<14359> A_IWL<14358> A_IWL<14357> A_IWL<14356> A_IWL<14355> A_IWL<14354> A_IWL<14353> A_IWL<14352> A_IWL<14351> A_IWL<14350> A_IWL<14349> A_IWL<14348> A_IWL<14347> A_IWL<14346> A_IWL<14345> A_IWL<14344> A_IWL<14343> A_IWL<14342> A_IWL<14341> A_IWL<14340> A_IWL<14339> A_IWL<14338> A_IWL<14337> A_IWL<14336> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<55> A_BLC<111> A_BLC<110> A_BLC_TOP<111> A_BLC_TOP<110> A_BLT<111> A_BLT<110> A_BLT_TOP<111> A_BLT_TOP<110> A_IWL<14079> A_IWL<14078> A_IWL<14077> A_IWL<14076> A_IWL<14075> A_IWL<14074> A_IWL<14073> A_IWL<14072> A_IWL<14071> A_IWL<14070> A_IWL<14069> A_IWL<14068> A_IWL<14067> A_IWL<14066> A_IWL<14065> A_IWL<14064> A_IWL<14063> A_IWL<14062> A_IWL<14061> A_IWL<14060> A_IWL<14059> A_IWL<14058> A_IWL<14057> A_IWL<14056> A_IWL<14055> A_IWL<14054> A_IWL<14053> A_IWL<14052> A_IWL<14051> A_IWL<14050> A_IWL<14049> A_IWL<14048> A_IWL<14047> A_IWL<14046> A_IWL<14045> A_IWL<14044> A_IWL<14043> A_IWL<14042> A_IWL<14041> A_IWL<14040> A_IWL<14039> A_IWL<14038> A_IWL<14037> A_IWL<14036> A_IWL<14035> A_IWL<14034> A_IWL<14033> A_IWL<14032> A_IWL<14031> A_IWL<14030> A_IWL<14029> A_IWL<14028> A_IWL<14027> A_IWL<14026> A_IWL<14025> A_IWL<14024> A_IWL<14023> A_IWL<14022> A_IWL<14021> A_IWL<14020> A_IWL<14019> A_IWL<14018> A_IWL<14017> A_IWL<14016> A_IWL<14015> A_IWL<14014> A_IWL<14013> A_IWL<14012> A_IWL<14011> A_IWL<14010> A_IWL<14009> A_IWL<14008> A_IWL<14007> A_IWL<14006> A_IWL<14005> A_IWL<14004> A_IWL<14003> A_IWL<14002> A_IWL<14001> A_IWL<14000> A_IWL<13999> A_IWL<13998> A_IWL<13997> A_IWL<13996> A_IWL<13995> A_IWL<13994> A_IWL<13993> A_IWL<13992> A_IWL<13991> A_IWL<13990> A_IWL<13989> A_IWL<13988> A_IWL<13987> A_IWL<13986> A_IWL<13985> A_IWL<13984> A_IWL<13983> A_IWL<13982> A_IWL<13981> A_IWL<13980> A_IWL<13979> A_IWL<13978> A_IWL<13977> A_IWL<13976> A_IWL<13975> A_IWL<13974> A_IWL<13973> A_IWL<13972> A_IWL<13971> A_IWL<13970> A_IWL<13969> A_IWL<13968> A_IWL<13967> A_IWL<13966> A_IWL<13965> A_IWL<13964> A_IWL<13963> A_IWL<13962> A_IWL<13961> A_IWL<13960> A_IWL<13959> A_IWL<13958> A_IWL<13957> A_IWL<13956> A_IWL<13955> A_IWL<13954> A_IWL<13953> A_IWL<13952> A_IWL<13951> A_IWL<13950> A_IWL<13949> A_IWL<13948> A_IWL<13947> A_IWL<13946> A_IWL<13945> A_IWL<13944> A_IWL<13943> A_IWL<13942> A_IWL<13941> A_IWL<13940> A_IWL<13939> A_IWL<13938> A_IWL<13937> A_IWL<13936> A_IWL<13935> A_IWL<13934> A_IWL<13933> A_IWL<13932> A_IWL<13931> A_IWL<13930> A_IWL<13929> A_IWL<13928> A_IWL<13927> A_IWL<13926> A_IWL<13925> A_IWL<13924> A_IWL<13923> A_IWL<13922> A_IWL<13921> A_IWL<13920> A_IWL<13919> A_IWL<13918> A_IWL<13917> A_IWL<13916> A_IWL<13915> A_IWL<13914> A_IWL<13913> A_IWL<13912> A_IWL<13911> A_IWL<13910> A_IWL<13909> A_IWL<13908> A_IWL<13907> A_IWL<13906> A_IWL<13905> A_IWL<13904> A_IWL<13903> A_IWL<13902> A_IWL<13901> A_IWL<13900> A_IWL<13899> A_IWL<13898> A_IWL<13897> A_IWL<13896> A_IWL<13895> A_IWL<13894> A_IWL<13893> A_IWL<13892> A_IWL<13891> A_IWL<13890> A_IWL<13889> A_IWL<13888> A_IWL<13887> A_IWL<13886> A_IWL<13885> A_IWL<13884> A_IWL<13883> A_IWL<13882> A_IWL<13881> A_IWL<13880> A_IWL<13879> A_IWL<13878> A_IWL<13877> A_IWL<13876> A_IWL<13875> A_IWL<13874> A_IWL<13873> A_IWL<13872> A_IWL<13871> A_IWL<13870> A_IWL<13869> A_IWL<13868> A_IWL<13867> A_IWL<13866> A_IWL<13865> A_IWL<13864> A_IWL<13863> A_IWL<13862> A_IWL<13861> A_IWL<13860> A_IWL<13859> A_IWL<13858> A_IWL<13857> A_IWL<13856> A_IWL<13855> A_IWL<13854> A_IWL<13853> A_IWL<13852> A_IWL<13851> A_IWL<13850> A_IWL<13849> A_IWL<13848> A_IWL<13847> A_IWL<13846> A_IWL<13845> A_IWL<13844> A_IWL<13843> A_IWL<13842> A_IWL<13841> A_IWL<13840> A_IWL<13839> A_IWL<13838> A_IWL<13837> A_IWL<13836> A_IWL<13835> A_IWL<13834> A_IWL<13833> A_IWL<13832> A_IWL<13831> A_IWL<13830> A_IWL<13829> A_IWL<13828> A_IWL<13827> A_IWL<13826> A_IWL<13825> A_IWL<13824> A_IWL<14335> A_IWL<14334> A_IWL<14333> A_IWL<14332> A_IWL<14331> A_IWL<14330> A_IWL<14329> A_IWL<14328> A_IWL<14327> A_IWL<14326> A_IWL<14325> A_IWL<14324> A_IWL<14323> A_IWL<14322> A_IWL<14321> A_IWL<14320> A_IWL<14319> A_IWL<14318> A_IWL<14317> A_IWL<14316> A_IWL<14315> A_IWL<14314> A_IWL<14313> A_IWL<14312> A_IWL<14311> A_IWL<14310> A_IWL<14309> A_IWL<14308> A_IWL<14307> A_IWL<14306> A_IWL<14305> A_IWL<14304> A_IWL<14303> A_IWL<14302> A_IWL<14301> A_IWL<14300> A_IWL<14299> A_IWL<14298> A_IWL<14297> A_IWL<14296> A_IWL<14295> A_IWL<14294> A_IWL<14293> A_IWL<14292> A_IWL<14291> A_IWL<14290> A_IWL<14289> A_IWL<14288> A_IWL<14287> A_IWL<14286> A_IWL<14285> A_IWL<14284> A_IWL<14283> A_IWL<14282> A_IWL<14281> A_IWL<14280> A_IWL<14279> A_IWL<14278> A_IWL<14277> A_IWL<14276> A_IWL<14275> A_IWL<14274> A_IWL<14273> A_IWL<14272> A_IWL<14271> A_IWL<14270> A_IWL<14269> A_IWL<14268> A_IWL<14267> A_IWL<14266> A_IWL<14265> A_IWL<14264> A_IWL<14263> A_IWL<14262> A_IWL<14261> A_IWL<14260> A_IWL<14259> A_IWL<14258> A_IWL<14257> A_IWL<14256> A_IWL<14255> A_IWL<14254> A_IWL<14253> A_IWL<14252> A_IWL<14251> A_IWL<14250> A_IWL<14249> A_IWL<14248> A_IWL<14247> A_IWL<14246> A_IWL<14245> A_IWL<14244> A_IWL<14243> A_IWL<14242> A_IWL<14241> A_IWL<14240> A_IWL<14239> A_IWL<14238> A_IWL<14237> A_IWL<14236> A_IWL<14235> A_IWL<14234> A_IWL<14233> A_IWL<14232> A_IWL<14231> A_IWL<14230> A_IWL<14229> A_IWL<14228> A_IWL<14227> A_IWL<14226> A_IWL<14225> A_IWL<14224> A_IWL<14223> A_IWL<14222> A_IWL<14221> A_IWL<14220> A_IWL<14219> A_IWL<14218> A_IWL<14217> A_IWL<14216> A_IWL<14215> A_IWL<14214> A_IWL<14213> A_IWL<14212> A_IWL<14211> A_IWL<14210> A_IWL<14209> A_IWL<14208> A_IWL<14207> A_IWL<14206> A_IWL<14205> A_IWL<14204> A_IWL<14203> A_IWL<14202> A_IWL<14201> A_IWL<14200> A_IWL<14199> A_IWL<14198> A_IWL<14197> A_IWL<14196> A_IWL<14195> A_IWL<14194> A_IWL<14193> A_IWL<14192> A_IWL<14191> A_IWL<14190> A_IWL<14189> A_IWL<14188> A_IWL<14187> A_IWL<14186> A_IWL<14185> A_IWL<14184> A_IWL<14183> A_IWL<14182> A_IWL<14181> A_IWL<14180> A_IWL<14179> A_IWL<14178> A_IWL<14177> A_IWL<14176> A_IWL<14175> A_IWL<14174> A_IWL<14173> A_IWL<14172> A_IWL<14171> A_IWL<14170> A_IWL<14169> A_IWL<14168> A_IWL<14167> A_IWL<14166> A_IWL<14165> A_IWL<14164> A_IWL<14163> A_IWL<14162> A_IWL<14161> A_IWL<14160> A_IWL<14159> A_IWL<14158> A_IWL<14157> A_IWL<14156> A_IWL<14155> A_IWL<14154> A_IWL<14153> A_IWL<14152> A_IWL<14151> A_IWL<14150> A_IWL<14149> A_IWL<14148> A_IWL<14147> A_IWL<14146> A_IWL<14145> A_IWL<14144> A_IWL<14143> A_IWL<14142> A_IWL<14141> A_IWL<14140> A_IWL<14139> A_IWL<14138> A_IWL<14137> A_IWL<14136> A_IWL<14135> A_IWL<14134> A_IWL<14133> A_IWL<14132> A_IWL<14131> A_IWL<14130> A_IWL<14129> A_IWL<14128> A_IWL<14127> A_IWL<14126> A_IWL<14125> A_IWL<14124> A_IWL<14123> A_IWL<14122> A_IWL<14121> A_IWL<14120> A_IWL<14119> A_IWL<14118> A_IWL<14117> A_IWL<14116> A_IWL<14115> A_IWL<14114> A_IWL<14113> A_IWL<14112> A_IWL<14111> A_IWL<14110> A_IWL<14109> A_IWL<14108> A_IWL<14107> A_IWL<14106> A_IWL<14105> A_IWL<14104> A_IWL<14103> A_IWL<14102> A_IWL<14101> A_IWL<14100> A_IWL<14099> A_IWL<14098> A_IWL<14097> A_IWL<14096> A_IWL<14095> A_IWL<14094> A_IWL<14093> A_IWL<14092> A_IWL<14091> A_IWL<14090> A_IWL<14089> A_IWL<14088> A_IWL<14087> A_IWL<14086> A_IWL<14085> A_IWL<14084> A_IWL<14083> A_IWL<14082> A_IWL<14081> A_IWL<14080> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<54> A_BLC<109> A_BLC<108> A_BLC_TOP<109> A_BLC_TOP<108> A_BLT<109> A_BLT<108> A_BLT_TOP<109> A_BLT_TOP<108> A_IWL<13823> A_IWL<13822> A_IWL<13821> A_IWL<13820> A_IWL<13819> A_IWL<13818> A_IWL<13817> A_IWL<13816> A_IWL<13815> A_IWL<13814> A_IWL<13813> A_IWL<13812> A_IWL<13811> A_IWL<13810> A_IWL<13809> A_IWL<13808> A_IWL<13807> A_IWL<13806> A_IWL<13805> A_IWL<13804> A_IWL<13803> A_IWL<13802> A_IWL<13801> A_IWL<13800> A_IWL<13799> A_IWL<13798> A_IWL<13797> A_IWL<13796> A_IWL<13795> A_IWL<13794> A_IWL<13793> A_IWL<13792> A_IWL<13791> A_IWL<13790> A_IWL<13789> A_IWL<13788> A_IWL<13787> A_IWL<13786> A_IWL<13785> A_IWL<13784> A_IWL<13783> A_IWL<13782> A_IWL<13781> A_IWL<13780> A_IWL<13779> A_IWL<13778> A_IWL<13777> A_IWL<13776> A_IWL<13775> A_IWL<13774> A_IWL<13773> A_IWL<13772> A_IWL<13771> A_IWL<13770> A_IWL<13769> A_IWL<13768> A_IWL<13767> A_IWL<13766> A_IWL<13765> A_IWL<13764> A_IWL<13763> A_IWL<13762> A_IWL<13761> A_IWL<13760> A_IWL<13759> A_IWL<13758> A_IWL<13757> A_IWL<13756> A_IWL<13755> A_IWL<13754> A_IWL<13753> A_IWL<13752> A_IWL<13751> A_IWL<13750> A_IWL<13749> A_IWL<13748> A_IWL<13747> A_IWL<13746> A_IWL<13745> A_IWL<13744> A_IWL<13743> A_IWL<13742> A_IWL<13741> A_IWL<13740> A_IWL<13739> A_IWL<13738> A_IWL<13737> A_IWL<13736> A_IWL<13735> A_IWL<13734> A_IWL<13733> A_IWL<13732> A_IWL<13731> A_IWL<13730> A_IWL<13729> A_IWL<13728> A_IWL<13727> A_IWL<13726> A_IWL<13725> A_IWL<13724> A_IWL<13723> A_IWL<13722> A_IWL<13721> A_IWL<13720> A_IWL<13719> A_IWL<13718> A_IWL<13717> A_IWL<13716> A_IWL<13715> A_IWL<13714> A_IWL<13713> A_IWL<13712> A_IWL<13711> A_IWL<13710> A_IWL<13709> A_IWL<13708> A_IWL<13707> A_IWL<13706> A_IWL<13705> A_IWL<13704> A_IWL<13703> A_IWL<13702> A_IWL<13701> A_IWL<13700> A_IWL<13699> A_IWL<13698> A_IWL<13697> A_IWL<13696> A_IWL<13695> A_IWL<13694> A_IWL<13693> A_IWL<13692> A_IWL<13691> A_IWL<13690> A_IWL<13689> A_IWL<13688> A_IWL<13687> A_IWL<13686> A_IWL<13685> A_IWL<13684> A_IWL<13683> A_IWL<13682> A_IWL<13681> A_IWL<13680> A_IWL<13679> A_IWL<13678> A_IWL<13677> A_IWL<13676> A_IWL<13675> A_IWL<13674> A_IWL<13673> A_IWL<13672> A_IWL<13671> A_IWL<13670> A_IWL<13669> A_IWL<13668> A_IWL<13667> A_IWL<13666> A_IWL<13665> A_IWL<13664> A_IWL<13663> A_IWL<13662> A_IWL<13661> A_IWL<13660> A_IWL<13659> A_IWL<13658> A_IWL<13657> A_IWL<13656> A_IWL<13655> A_IWL<13654> A_IWL<13653> A_IWL<13652> A_IWL<13651> A_IWL<13650> A_IWL<13649> A_IWL<13648> A_IWL<13647> A_IWL<13646> A_IWL<13645> A_IWL<13644> A_IWL<13643> A_IWL<13642> A_IWL<13641> A_IWL<13640> A_IWL<13639> A_IWL<13638> A_IWL<13637> A_IWL<13636> A_IWL<13635> A_IWL<13634> A_IWL<13633> A_IWL<13632> A_IWL<13631> A_IWL<13630> A_IWL<13629> A_IWL<13628> A_IWL<13627> A_IWL<13626> A_IWL<13625> A_IWL<13624> A_IWL<13623> A_IWL<13622> A_IWL<13621> A_IWL<13620> A_IWL<13619> A_IWL<13618> A_IWL<13617> A_IWL<13616> A_IWL<13615> A_IWL<13614> A_IWL<13613> A_IWL<13612> A_IWL<13611> A_IWL<13610> A_IWL<13609> A_IWL<13608> A_IWL<13607> A_IWL<13606> A_IWL<13605> A_IWL<13604> A_IWL<13603> A_IWL<13602> A_IWL<13601> A_IWL<13600> A_IWL<13599> A_IWL<13598> A_IWL<13597> A_IWL<13596> A_IWL<13595> A_IWL<13594> A_IWL<13593> A_IWL<13592> A_IWL<13591> A_IWL<13590> A_IWL<13589> A_IWL<13588> A_IWL<13587> A_IWL<13586> A_IWL<13585> A_IWL<13584> A_IWL<13583> A_IWL<13582> A_IWL<13581> A_IWL<13580> A_IWL<13579> A_IWL<13578> A_IWL<13577> A_IWL<13576> A_IWL<13575> A_IWL<13574> A_IWL<13573> A_IWL<13572> A_IWL<13571> A_IWL<13570> A_IWL<13569> A_IWL<13568> A_IWL<14079> A_IWL<14078> A_IWL<14077> A_IWL<14076> A_IWL<14075> A_IWL<14074> A_IWL<14073> A_IWL<14072> A_IWL<14071> A_IWL<14070> A_IWL<14069> A_IWL<14068> A_IWL<14067> A_IWL<14066> A_IWL<14065> A_IWL<14064> A_IWL<14063> A_IWL<14062> A_IWL<14061> A_IWL<14060> A_IWL<14059> A_IWL<14058> A_IWL<14057> A_IWL<14056> A_IWL<14055> A_IWL<14054> A_IWL<14053> A_IWL<14052> A_IWL<14051> A_IWL<14050> A_IWL<14049> A_IWL<14048> A_IWL<14047> A_IWL<14046> A_IWL<14045> A_IWL<14044> A_IWL<14043> A_IWL<14042> A_IWL<14041> A_IWL<14040> A_IWL<14039> A_IWL<14038> A_IWL<14037> A_IWL<14036> A_IWL<14035> A_IWL<14034> A_IWL<14033> A_IWL<14032> A_IWL<14031> A_IWL<14030> A_IWL<14029> A_IWL<14028> A_IWL<14027> A_IWL<14026> A_IWL<14025> A_IWL<14024> A_IWL<14023> A_IWL<14022> A_IWL<14021> A_IWL<14020> A_IWL<14019> A_IWL<14018> A_IWL<14017> A_IWL<14016> A_IWL<14015> A_IWL<14014> A_IWL<14013> A_IWL<14012> A_IWL<14011> A_IWL<14010> A_IWL<14009> A_IWL<14008> A_IWL<14007> A_IWL<14006> A_IWL<14005> A_IWL<14004> A_IWL<14003> A_IWL<14002> A_IWL<14001> A_IWL<14000> A_IWL<13999> A_IWL<13998> A_IWL<13997> A_IWL<13996> A_IWL<13995> A_IWL<13994> A_IWL<13993> A_IWL<13992> A_IWL<13991> A_IWL<13990> A_IWL<13989> A_IWL<13988> A_IWL<13987> A_IWL<13986> A_IWL<13985> A_IWL<13984> A_IWL<13983> A_IWL<13982> A_IWL<13981> A_IWL<13980> A_IWL<13979> A_IWL<13978> A_IWL<13977> A_IWL<13976> A_IWL<13975> A_IWL<13974> A_IWL<13973> A_IWL<13972> A_IWL<13971> A_IWL<13970> A_IWL<13969> A_IWL<13968> A_IWL<13967> A_IWL<13966> A_IWL<13965> A_IWL<13964> A_IWL<13963> A_IWL<13962> A_IWL<13961> A_IWL<13960> A_IWL<13959> A_IWL<13958> A_IWL<13957> A_IWL<13956> A_IWL<13955> A_IWL<13954> A_IWL<13953> A_IWL<13952> A_IWL<13951> A_IWL<13950> A_IWL<13949> A_IWL<13948> A_IWL<13947> A_IWL<13946> A_IWL<13945> A_IWL<13944> A_IWL<13943> A_IWL<13942> A_IWL<13941> A_IWL<13940> A_IWL<13939> A_IWL<13938> A_IWL<13937> A_IWL<13936> A_IWL<13935> A_IWL<13934> A_IWL<13933> A_IWL<13932> A_IWL<13931> A_IWL<13930> A_IWL<13929> A_IWL<13928> A_IWL<13927> A_IWL<13926> A_IWL<13925> A_IWL<13924> A_IWL<13923> A_IWL<13922> A_IWL<13921> A_IWL<13920> A_IWL<13919> A_IWL<13918> A_IWL<13917> A_IWL<13916> A_IWL<13915> A_IWL<13914> A_IWL<13913> A_IWL<13912> A_IWL<13911> A_IWL<13910> A_IWL<13909> A_IWL<13908> A_IWL<13907> A_IWL<13906> A_IWL<13905> A_IWL<13904> A_IWL<13903> A_IWL<13902> A_IWL<13901> A_IWL<13900> A_IWL<13899> A_IWL<13898> A_IWL<13897> A_IWL<13896> A_IWL<13895> A_IWL<13894> A_IWL<13893> A_IWL<13892> A_IWL<13891> A_IWL<13890> A_IWL<13889> A_IWL<13888> A_IWL<13887> A_IWL<13886> A_IWL<13885> A_IWL<13884> A_IWL<13883> A_IWL<13882> A_IWL<13881> A_IWL<13880> A_IWL<13879> A_IWL<13878> A_IWL<13877> A_IWL<13876> A_IWL<13875> A_IWL<13874> A_IWL<13873> A_IWL<13872> A_IWL<13871> A_IWL<13870> A_IWL<13869> A_IWL<13868> A_IWL<13867> A_IWL<13866> A_IWL<13865> A_IWL<13864> A_IWL<13863> A_IWL<13862> A_IWL<13861> A_IWL<13860> A_IWL<13859> A_IWL<13858> A_IWL<13857> A_IWL<13856> A_IWL<13855> A_IWL<13854> A_IWL<13853> A_IWL<13852> A_IWL<13851> A_IWL<13850> A_IWL<13849> A_IWL<13848> A_IWL<13847> A_IWL<13846> A_IWL<13845> A_IWL<13844> A_IWL<13843> A_IWL<13842> A_IWL<13841> A_IWL<13840> A_IWL<13839> A_IWL<13838> A_IWL<13837> A_IWL<13836> A_IWL<13835> A_IWL<13834> A_IWL<13833> A_IWL<13832> A_IWL<13831> A_IWL<13830> A_IWL<13829> A_IWL<13828> A_IWL<13827> A_IWL<13826> A_IWL<13825> A_IWL<13824> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<53> A_BLC<107> A_BLC<106> A_BLC_TOP<107> A_BLC_TOP<106> A_BLT<107> A_BLT<106> A_BLT_TOP<107> A_BLT_TOP<106> A_IWL<13567> A_IWL<13566> A_IWL<13565> A_IWL<13564> A_IWL<13563> A_IWL<13562> A_IWL<13561> A_IWL<13560> A_IWL<13559> A_IWL<13558> A_IWL<13557> A_IWL<13556> A_IWL<13555> A_IWL<13554> A_IWL<13553> A_IWL<13552> A_IWL<13551> A_IWL<13550> A_IWL<13549> A_IWL<13548> A_IWL<13547> A_IWL<13546> A_IWL<13545> A_IWL<13544> A_IWL<13543> A_IWL<13542> A_IWL<13541> A_IWL<13540> A_IWL<13539> A_IWL<13538> A_IWL<13537> A_IWL<13536> A_IWL<13535> A_IWL<13534> A_IWL<13533> A_IWL<13532> A_IWL<13531> A_IWL<13530> A_IWL<13529> A_IWL<13528> A_IWL<13527> A_IWL<13526> A_IWL<13525> A_IWL<13524> A_IWL<13523> A_IWL<13522> A_IWL<13521> A_IWL<13520> A_IWL<13519> A_IWL<13518> A_IWL<13517> A_IWL<13516> A_IWL<13515> A_IWL<13514> A_IWL<13513> A_IWL<13512> A_IWL<13511> A_IWL<13510> A_IWL<13509> A_IWL<13508> A_IWL<13507> A_IWL<13506> A_IWL<13505> A_IWL<13504> A_IWL<13503> A_IWL<13502> A_IWL<13501> A_IWL<13500> A_IWL<13499> A_IWL<13498> A_IWL<13497> A_IWL<13496> A_IWL<13495> A_IWL<13494> A_IWL<13493> A_IWL<13492> A_IWL<13491> A_IWL<13490> A_IWL<13489> A_IWL<13488> A_IWL<13487> A_IWL<13486> A_IWL<13485> A_IWL<13484> A_IWL<13483> A_IWL<13482> A_IWL<13481> A_IWL<13480> A_IWL<13479> A_IWL<13478> A_IWL<13477> A_IWL<13476> A_IWL<13475> A_IWL<13474> A_IWL<13473> A_IWL<13472> A_IWL<13471> A_IWL<13470> A_IWL<13469> A_IWL<13468> A_IWL<13467> A_IWL<13466> A_IWL<13465> A_IWL<13464> A_IWL<13463> A_IWL<13462> A_IWL<13461> A_IWL<13460> A_IWL<13459> A_IWL<13458> A_IWL<13457> A_IWL<13456> A_IWL<13455> A_IWL<13454> A_IWL<13453> A_IWL<13452> A_IWL<13451> A_IWL<13450> A_IWL<13449> A_IWL<13448> A_IWL<13447> A_IWL<13446> A_IWL<13445> A_IWL<13444> A_IWL<13443> A_IWL<13442> A_IWL<13441> A_IWL<13440> A_IWL<13439> A_IWL<13438> A_IWL<13437> A_IWL<13436> A_IWL<13435> A_IWL<13434> A_IWL<13433> A_IWL<13432> A_IWL<13431> A_IWL<13430> A_IWL<13429> A_IWL<13428> A_IWL<13427> A_IWL<13426> A_IWL<13425> A_IWL<13424> A_IWL<13423> A_IWL<13422> A_IWL<13421> A_IWL<13420> A_IWL<13419> A_IWL<13418> A_IWL<13417> A_IWL<13416> A_IWL<13415> A_IWL<13414> A_IWL<13413> A_IWL<13412> A_IWL<13411> A_IWL<13410> A_IWL<13409> A_IWL<13408> A_IWL<13407> A_IWL<13406> A_IWL<13405> A_IWL<13404> A_IWL<13403> A_IWL<13402> A_IWL<13401> A_IWL<13400> A_IWL<13399> A_IWL<13398> A_IWL<13397> A_IWL<13396> A_IWL<13395> A_IWL<13394> A_IWL<13393> A_IWL<13392> A_IWL<13391> A_IWL<13390> A_IWL<13389> A_IWL<13388> A_IWL<13387> A_IWL<13386> A_IWL<13385> A_IWL<13384> A_IWL<13383> A_IWL<13382> A_IWL<13381> A_IWL<13380> A_IWL<13379> A_IWL<13378> A_IWL<13377> A_IWL<13376> A_IWL<13375> A_IWL<13374> A_IWL<13373> A_IWL<13372> A_IWL<13371> A_IWL<13370> A_IWL<13369> A_IWL<13368> A_IWL<13367> A_IWL<13366> A_IWL<13365> A_IWL<13364> A_IWL<13363> A_IWL<13362> A_IWL<13361> A_IWL<13360> A_IWL<13359> A_IWL<13358> A_IWL<13357> A_IWL<13356> A_IWL<13355> A_IWL<13354> A_IWL<13353> A_IWL<13352> A_IWL<13351> A_IWL<13350> A_IWL<13349> A_IWL<13348> A_IWL<13347> A_IWL<13346> A_IWL<13345> A_IWL<13344> A_IWL<13343> A_IWL<13342> A_IWL<13341> A_IWL<13340> A_IWL<13339> A_IWL<13338> A_IWL<13337> A_IWL<13336> A_IWL<13335> A_IWL<13334> A_IWL<13333> A_IWL<13332> A_IWL<13331> A_IWL<13330> A_IWL<13329> A_IWL<13328> A_IWL<13327> A_IWL<13326> A_IWL<13325> A_IWL<13324> A_IWL<13323> A_IWL<13322> A_IWL<13321> A_IWL<13320> A_IWL<13319> A_IWL<13318> A_IWL<13317> A_IWL<13316> A_IWL<13315> A_IWL<13314> A_IWL<13313> A_IWL<13312> A_IWL<13823> A_IWL<13822> A_IWL<13821> A_IWL<13820> A_IWL<13819> A_IWL<13818> A_IWL<13817> A_IWL<13816> A_IWL<13815> A_IWL<13814> A_IWL<13813> A_IWL<13812> A_IWL<13811> A_IWL<13810> A_IWL<13809> A_IWL<13808> A_IWL<13807> A_IWL<13806> A_IWL<13805> A_IWL<13804> A_IWL<13803> A_IWL<13802> A_IWL<13801> A_IWL<13800> A_IWL<13799> A_IWL<13798> A_IWL<13797> A_IWL<13796> A_IWL<13795> A_IWL<13794> A_IWL<13793> A_IWL<13792> A_IWL<13791> A_IWL<13790> A_IWL<13789> A_IWL<13788> A_IWL<13787> A_IWL<13786> A_IWL<13785> A_IWL<13784> A_IWL<13783> A_IWL<13782> A_IWL<13781> A_IWL<13780> A_IWL<13779> A_IWL<13778> A_IWL<13777> A_IWL<13776> A_IWL<13775> A_IWL<13774> A_IWL<13773> A_IWL<13772> A_IWL<13771> A_IWL<13770> A_IWL<13769> A_IWL<13768> A_IWL<13767> A_IWL<13766> A_IWL<13765> A_IWL<13764> A_IWL<13763> A_IWL<13762> A_IWL<13761> A_IWL<13760> A_IWL<13759> A_IWL<13758> A_IWL<13757> A_IWL<13756> A_IWL<13755> A_IWL<13754> A_IWL<13753> A_IWL<13752> A_IWL<13751> A_IWL<13750> A_IWL<13749> A_IWL<13748> A_IWL<13747> A_IWL<13746> A_IWL<13745> A_IWL<13744> A_IWL<13743> A_IWL<13742> A_IWL<13741> A_IWL<13740> A_IWL<13739> A_IWL<13738> A_IWL<13737> A_IWL<13736> A_IWL<13735> A_IWL<13734> A_IWL<13733> A_IWL<13732> A_IWL<13731> A_IWL<13730> A_IWL<13729> A_IWL<13728> A_IWL<13727> A_IWL<13726> A_IWL<13725> A_IWL<13724> A_IWL<13723> A_IWL<13722> A_IWL<13721> A_IWL<13720> A_IWL<13719> A_IWL<13718> A_IWL<13717> A_IWL<13716> A_IWL<13715> A_IWL<13714> A_IWL<13713> A_IWL<13712> A_IWL<13711> A_IWL<13710> A_IWL<13709> A_IWL<13708> A_IWL<13707> A_IWL<13706> A_IWL<13705> A_IWL<13704> A_IWL<13703> A_IWL<13702> A_IWL<13701> A_IWL<13700> A_IWL<13699> A_IWL<13698> A_IWL<13697> A_IWL<13696> A_IWL<13695> A_IWL<13694> A_IWL<13693> A_IWL<13692> A_IWL<13691> A_IWL<13690> A_IWL<13689> A_IWL<13688> A_IWL<13687> A_IWL<13686> A_IWL<13685> A_IWL<13684> A_IWL<13683> A_IWL<13682> A_IWL<13681> A_IWL<13680> A_IWL<13679> A_IWL<13678> A_IWL<13677> A_IWL<13676> A_IWL<13675> A_IWL<13674> A_IWL<13673> A_IWL<13672> A_IWL<13671> A_IWL<13670> A_IWL<13669> A_IWL<13668> A_IWL<13667> A_IWL<13666> A_IWL<13665> A_IWL<13664> A_IWL<13663> A_IWL<13662> A_IWL<13661> A_IWL<13660> A_IWL<13659> A_IWL<13658> A_IWL<13657> A_IWL<13656> A_IWL<13655> A_IWL<13654> A_IWL<13653> A_IWL<13652> A_IWL<13651> A_IWL<13650> A_IWL<13649> A_IWL<13648> A_IWL<13647> A_IWL<13646> A_IWL<13645> A_IWL<13644> A_IWL<13643> A_IWL<13642> A_IWL<13641> A_IWL<13640> A_IWL<13639> A_IWL<13638> A_IWL<13637> A_IWL<13636> A_IWL<13635> A_IWL<13634> A_IWL<13633> A_IWL<13632> A_IWL<13631> A_IWL<13630> A_IWL<13629> A_IWL<13628> A_IWL<13627> A_IWL<13626> A_IWL<13625> A_IWL<13624> A_IWL<13623> A_IWL<13622> A_IWL<13621> A_IWL<13620> A_IWL<13619> A_IWL<13618> A_IWL<13617> A_IWL<13616> A_IWL<13615> A_IWL<13614> A_IWL<13613> A_IWL<13612> A_IWL<13611> A_IWL<13610> A_IWL<13609> A_IWL<13608> A_IWL<13607> A_IWL<13606> A_IWL<13605> A_IWL<13604> A_IWL<13603> A_IWL<13602> A_IWL<13601> A_IWL<13600> A_IWL<13599> A_IWL<13598> A_IWL<13597> A_IWL<13596> A_IWL<13595> A_IWL<13594> A_IWL<13593> A_IWL<13592> A_IWL<13591> A_IWL<13590> A_IWL<13589> A_IWL<13588> A_IWL<13587> A_IWL<13586> A_IWL<13585> A_IWL<13584> A_IWL<13583> A_IWL<13582> A_IWL<13581> A_IWL<13580> A_IWL<13579> A_IWL<13578> A_IWL<13577> A_IWL<13576> A_IWL<13575> A_IWL<13574> A_IWL<13573> A_IWL<13572> A_IWL<13571> A_IWL<13570> A_IWL<13569> A_IWL<13568> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<52> A_BLC<105> A_BLC<104> A_BLC_TOP<105> A_BLC_TOP<104> A_BLT<105> A_BLT<104> A_BLT_TOP<105> A_BLT_TOP<104> A_IWL<13311> A_IWL<13310> A_IWL<13309> A_IWL<13308> A_IWL<13307> A_IWL<13306> A_IWL<13305> A_IWL<13304> A_IWL<13303> A_IWL<13302> A_IWL<13301> A_IWL<13300> A_IWL<13299> A_IWL<13298> A_IWL<13297> A_IWL<13296> A_IWL<13295> A_IWL<13294> A_IWL<13293> A_IWL<13292> A_IWL<13291> A_IWL<13290> A_IWL<13289> A_IWL<13288> A_IWL<13287> A_IWL<13286> A_IWL<13285> A_IWL<13284> A_IWL<13283> A_IWL<13282> A_IWL<13281> A_IWL<13280> A_IWL<13279> A_IWL<13278> A_IWL<13277> A_IWL<13276> A_IWL<13275> A_IWL<13274> A_IWL<13273> A_IWL<13272> A_IWL<13271> A_IWL<13270> A_IWL<13269> A_IWL<13268> A_IWL<13267> A_IWL<13266> A_IWL<13265> A_IWL<13264> A_IWL<13263> A_IWL<13262> A_IWL<13261> A_IWL<13260> A_IWL<13259> A_IWL<13258> A_IWL<13257> A_IWL<13256> A_IWL<13255> A_IWL<13254> A_IWL<13253> A_IWL<13252> A_IWL<13251> A_IWL<13250> A_IWL<13249> A_IWL<13248> A_IWL<13247> A_IWL<13246> A_IWL<13245> A_IWL<13244> A_IWL<13243> A_IWL<13242> A_IWL<13241> A_IWL<13240> A_IWL<13239> A_IWL<13238> A_IWL<13237> A_IWL<13236> A_IWL<13235> A_IWL<13234> A_IWL<13233> A_IWL<13232> A_IWL<13231> A_IWL<13230> A_IWL<13229> A_IWL<13228> A_IWL<13227> A_IWL<13226> A_IWL<13225> A_IWL<13224> A_IWL<13223> A_IWL<13222> A_IWL<13221> A_IWL<13220> A_IWL<13219> A_IWL<13218> A_IWL<13217> A_IWL<13216> A_IWL<13215> A_IWL<13214> A_IWL<13213> A_IWL<13212> A_IWL<13211> A_IWL<13210> A_IWL<13209> A_IWL<13208> A_IWL<13207> A_IWL<13206> A_IWL<13205> A_IWL<13204> A_IWL<13203> A_IWL<13202> A_IWL<13201> A_IWL<13200> A_IWL<13199> A_IWL<13198> A_IWL<13197> A_IWL<13196> A_IWL<13195> A_IWL<13194> A_IWL<13193> A_IWL<13192> A_IWL<13191> A_IWL<13190> A_IWL<13189> A_IWL<13188> A_IWL<13187> A_IWL<13186> A_IWL<13185> A_IWL<13184> A_IWL<13183> A_IWL<13182> A_IWL<13181> A_IWL<13180> A_IWL<13179> A_IWL<13178> A_IWL<13177> A_IWL<13176> A_IWL<13175> A_IWL<13174> A_IWL<13173> A_IWL<13172> A_IWL<13171> A_IWL<13170> A_IWL<13169> A_IWL<13168> A_IWL<13167> A_IWL<13166> A_IWL<13165> A_IWL<13164> A_IWL<13163> A_IWL<13162> A_IWL<13161> A_IWL<13160> A_IWL<13159> A_IWL<13158> A_IWL<13157> A_IWL<13156> A_IWL<13155> A_IWL<13154> A_IWL<13153> A_IWL<13152> A_IWL<13151> A_IWL<13150> A_IWL<13149> A_IWL<13148> A_IWL<13147> A_IWL<13146> A_IWL<13145> A_IWL<13144> A_IWL<13143> A_IWL<13142> A_IWL<13141> A_IWL<13140> A_IWL<13139> A_IWL<13138> A_IWL<13137> A_IWL<13136> A_IWL<13135> A_IWL<13134> A_IWL<13133> A_IWL<13132> A_IWL<13131> A_IWL<13130> A_IWL<13129> A_IWL<13128> A_IWL<13127> A_IWL<13126> A_IWL<13125> A_IWL<13124> A_IWL<13123> A_IWL<13122> A_IWL<13121> A_IWL<13120> A_IWL<13119> A_IWL<13118> A_IWL<13117> A_IWL<13116> A_IWL<13115> A_IWL<13114> A_IWL<13113> A_IWL<13112> A_IWL<13111> A_IWL<13110> A_IWL<13109> A_IWL<13108> A_IWL<13107> A_IWL<13106> A_IWL<13105> A_IWL<13104> A_IWL<13103> A_IWL<13102> A_IWL<13101> A_IWL<13100> A_IWL<13099> A_IWL<13098> A_IWL<13097> A_IWL<13096> A_IWL<13095> A_IWL<13094> A_IWL<13093> A_IWL<13092> A_IWL<13091> A_IWL<13090> A_IWL<13089> A_IWL<13088> A_IWL<13087> A_IWL<13086> A_IWL<13085> A_IWL<13084> A_IWL<13083> A_IWL<13082> A_IWL<13081> A_IWL<13080> A_IWL<13079> A_IWL<13078> A_IWL<13077> A_IWL<13076> A_IWL<13075> A_IWL<13074> A_IWL<13073> A_IWL<13072> A_IWL<13071> A_IWL<13070> A_IWL<13069> A_IWL<13068> A_IWL<13067> A_IWL<13066> A_IWL<13065> A_IWL<13064> A_IWL<13063> A_IWL<13062> A_IWL<13061> A_IWL<13060> A_IWL<13059> A_IWL<13058> A_IWL<13057> A_IWL<13056> A_IWL<13567> A_IWL<13566> A_IWL<13565> A_IWL<13564> A_IWL<13563> A_IWL<13562> A_IWL<13561> A_IWL<13560> A_IWL<13559> A_IWL<13558> A_IWL<13557> A_IWL<13556> A_IWL<13555> A_IWL<13554> A_IWL<13553> A_IWL<13552> A_IWL<13551> A_IWL<13550> A_IWL<13549> A_IWL<13548> A_IWL<13547> A_IWL<13546> A_IWL<13545> A_IWL<13544> A_IWL<13543> A_IWL<13542> A_IWL<13541> A_IWL<13540> A_IWL<13539> A_IWL<13538> A_IWL<13537> A_IWL<13536> A_IWL<13535> A_IWL<13534> A_IWL<13533> A_IWL<13532> A_IWL<13531> A_IWL<13530> A_IWL<13529> A_IWL<13528> A_IWL<13527> A_IWL<13526> A_IWL<13525> A_IWL<13524> A_IWL<13523> A_IWL<13522> A_IWL<13521> A_IWL<13520> A_IWL<13519> A_IWL<13518> A_IWL<13517> A_IWL<13516> A_IWL<13515> A_IWL<13514> A_IWL<13513> A_IWL<13512> A_IWL<13511> A_IWL<13510> A_IWL<13509> A_IWL<13508> A_IWL<13507> A_IWL<13506> A_IWL<13505> A_IWL<13504> A_IWL<13503> A_IWL<13502> A_IWL<13501> A_IWL<13500> A_IWL<13499> A_IWL<13498> A_IWL<13497> A_IWL<13496> A_IWL<13495> A_IWL<13494> A_IWL<13493> A_IWL<13492> A_IWL<13491> A_IWL<13490> A_IWL<13489> A_IWL<13488> A_IWL<13487> A_IWL<13486> A_IWL<13485> A_IWL<13484> A_IWL<13483> A_IWL<13482> A_IWL<13481> A_IWL<13480> A_IWL<13479> A_IWL<13478> A_IWL<13477> A_IWL<13476> A_IWL<13475> A_IWL<13474> A_IWL<13473> A_IWL<13472> A_IWL<13471> A_IWL<13470> A_IWL<13469> A_IWL<13468> A_IWL<13467> A_IWL<13466> A_IWL<13465> A_IWL<13464> A_IWL<13463> A_IWL<13462> A_IWL<13461> A_IWL<13460> A_IWL<13459> A_IWL<13458> A_IWL<13457> A_IWL<13456> A_IWL<13455> A_IWL<13454> A_IWL<13453> A_IWL<13452> A_IWL<13451> A_IWL<13450> A_IWL<13449> A_IWL<13448> A_IWL<13447> A_IWL<13446> A_IWL<13445> A_IWL<13444> A_IWL<13443> A_IWL<13442> A_IWL<13441> A_IWL<13440> A_IWL<13439> A_IWL<13438> A_IWL<13437> A_IWL<13436> A_IWL<13435> A_IWL<13434> A_IWL<13433> A_IWL<13432> A_IWL<13431> A_IWL<13430> A_IWL<13429> A_IWL<13428> A_IWL<13427> A_IWL<13426> A_IWL<13425> A_IWL<13424> A_IWL<13423> A_IWL<13422> A_IWL<13421> A_IWL<13420> A_IWL<13419> A_IWL<13418> A_IWL<13417> A_IWL<13416> A_IWL<13415> A_IWL<13414> A_IWL<13413> A_IWL<13412> A_IWL<13411> A_IWL<13410> A_IWL<13409> A_IWL<13408> A_IWL<13407> A_IWL<13406> A_IWL<13405> A_IWL<13404> A_IWL<13403> A_IWL<13402> A_IWL<13401> A_IWL<13400> A_IWL<13399> A_IWL<13398> A_IWL<13397> A_IWL<13396> A_IWL<13395> A_IWL<13394> A_IWL<13393> A_IWL<13392> A_IWL<13391> A_IWL<13390> A_IWL<13389> A_IWL<13388> A_IWL<13387> A_IWL<13386> A_IWL<13385> A_IWL<13384> A_IWL<13383> A_IWL<13382> A_IWL<13381> A_IWL<13380> A_IWL<13379> A_IWL<13378> A_IWL<13377> A_IWL<13376> A_IWL<13375> A_IWL<13374> A_IWL<13373> A_IWL<13372> A_IWL<13371> A_IWL<13370> A_IWL<13369> A_IWL<13368> A_IWL<13367> A_IWL<13366> A_IWL<13365> A_IWL<13364> A_IWL<13363> A_IWL<13362> A_IWL<13361> A_IWL<13360> A_IWL<13359> A_IWL<13358> A_IWL<13357> A_IWL<13356> A_IWL<13355> A_IWL<13354> A_IWL<13353> A_IWL<13352> A_IWL<13351> A_IWL<13350> A_IWL<13349> A_IWL<13348> A_IWL<13347> A_IWL<13346> A_IWL<13345> A_IWL<13344> A_IWL<13343> A_IWL<13342> A_IWL<13341> A_IWL<13340> A_IWL<13339> A_IWL<13338> A_IWL<13337> A_IWL<13336> A_IWL<13335> A_IWL<13334> A_IWL<13333> A_IWL<13332> A_IWL<13331> A_IWL<13330> A_IWL<13329> A_IWL<13328> A_IWL<13327> A_IWL<13326> A_IWL<13325> A_IWL<13324> A_IWL<13323> A_IWL<13322> A_IWL<13321> A_IWL<13320> A_IWL<13319> A_IWL<13318> A_IWL<13317> A_IWL<13316> A_IWL<13315> A_IWL<13314> A_IWL<13313> A_IWL<13312> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<51> A_BLC<103> A_BLC<102> A_BLC_TOP<103> A_BLC_TOP<102> A_BLT<103> A_BLT<102> A_BLT_TOP<103> A_BLT_TOP<102> A_IWL<13055> A_IWL<13054> A_IWL<13053> A_IWL<13052> A_IWL<13051> A_IWL<13050> A_IWL<13049> A_IWL<13048> A_IWL<13047> A_IWL<13046> A_IWL<13045> A_IWL<13044> A_IWL<13043> A_IWL<13042> A_IWL<13041> A_IWL<13040> A_IWL<13039> A_IWL<13038> A_IWL<13037> A_IWL<13036> A_IWL<13035> A_IWL<13034> A_IWL<13033> A_IWL<13032> A_IWL<13031> A_IWL<13030> A_IWL<13029> A_IWL<13028> A_IWL<13027> A_IWL<13026> A_IWL<13025> A_IWL<13024> A_IWL<13023> A_IWL<13022> A_IWL<13021> A_IWL<13020> A_IWL<13019> A_IWL<13018> A_IWL<13017> A_IWL<13016> A_IWL<13015> A_IWL<13014> A_IWL<13013> A_IWL<13012> A_IWL<13011> A_IWL<13010> A_IWL<13009> A_IWL<13008> A_IWL<13007> A_IWL<13006> A_IWL<13005> A_IWL<13004> A_IWL<13003> A_IWL<13002> A_IWL<13001> A_IWL<13000> A_IWL<12999> A_IWL<12998> A_IWL<12997> A_IWL<12996> A_IWL<12995> A_IWL<12994> A_IWL<12993> A_IWL<12992> A_IWL<12991> A_IWL<12990> A_IWL<12989> A_IWL<12988> A_IWL<12987> A_IWL<12986> A_IWL<12985> A_IWL<12984> A_IWL<12983> A_IWL<12982> A_IWL<12981> A_IWL<12980> A_IWL<12979> A_IWL<12978> A_IWL<12977> A_IWL<12976> A_IWL<12975> A_IWL<12974> A_IWL<12973> A_IWL<12972> A_IWL<12971> A_IWL<12970> A_IWL<12969> A_IWL<12968> A_IWL<12967> A_IWL<12966> A_IWL<12965> A_IWL<12964> A_IWL<12963> A_IWL<12962> A_IWL<12961> A_IWL<12960> A_IWL<12959> A_IWL<12958> A_IWL<12957> A_IWL<12956> A_IWL<12955> A_IWL<12954> A_IWL<12953> A_IWL<12952> A_IWL<12951> A_IWL<12950> A_IWL<12949> A_IWL<12948> A_IWL<12947> A_IWL<12946> A_IWL<12945> A_IWL<12944> A_IWL<12943> A_IWL<12942> A_IWL<12941> A_IWL<12940> A_IWL<12939> A_IWL<12938> A_IWL<12937> A_IWL<12936> A_IWL<12935> A_IWL<12934> A_IWL<12933> A_IWL<12932> A_IWL<12931> A_IWL<12930> A_IWL<12929> A_IWL<12928> A_IWL<12927> A_IWL<12926> A_IWL<12925> A_IWL<12924> A_IWL<12923> A_IWL<12922> A_IWL<12921> A_IWL<12920> A_IWL<12919> A_IWL<12918> A_IWL<12917> A_IWL<12916> A_IWL<12915> A_IWL<12914> A_IWL<12913> A_IWL<12912> A_IWL<12911> A_IWL<12910> A_IWL<12909> A_IWL<12908> A_IWL<12907> A_IWL<12906> A_IWL<12905> A_IWL<12904> A_IWL<12903> A_IWL<12902> A_IWL<12901> A_IWL<12900> A_IWL<12899> A_IWL<12898> A_IWL<12897> A_IWL<12896> A_IWL<12895> A_IWL<12894> A_IWL<12893> A_IWL<12892> A_IWL<12891> A_IWL<12890> A_IWL<12889> A_IWL<12888> A_IWL<12887> A_IWL<12886> A_IWL<12885> A_IWL<12884> A_IWL<12883> A_IWL<12882> A_IWL<12881> A_IWL<12880> A_IWL<12879> A_IWL<12878> A_IWL<12877> A_IWL<12876> A_IWL<12875> A_IWL<12874> A_IWL<12873> A_IWL<12872> A_IWL<12871> A_IWL<12870> A_IWL<12869> A_IWL<12868> A_IWL<12867> A_IWL<12866> A_IWL<12865> A_IWL<12864> A_IWL<12863> A_IWL<12862> A_IWL<12861> A_IWL<12860> A_IWL<12859> A_IWL<12858> A_IWL<12857> A_IWL<12856> A_IWL<12855> A_IWL<12854> A_IWL<12853> A_IWL<12852> A_IWL<12851> A_IWL<12850> A_IWL<12849> A_IWL<12848> A_IWL<12847> A_IWL<12846> A_IWL<12845> A_IWL<12844> A_IWL<12843> A_IWL<12842> A_IWL<12841> A_IWL<12840> A_IWL<12839> A_IWL<12838> A_IWL<12837> A_IWL<12836> A_IWL<12835> A_IWL<12834> A_IWL<12833> A_IWL<12832> A_IWL<12831> A_IWL<12830> A_IWL<12829> A_IWL<12828> A_IWL<12827> A_IWL<12826> A_IWL<12825> A_IWL<12824> A_IWL<12823> A_IWL<12822> A_IWL<12821> A_IWL<12820> A_IWL<12819> A_IWL<12818> A_IWL<12817> A_IWL<12816> A_IWL<12815> A_IWL<12814> A_IWL<12813> A_IWL<12812> A_IWL<12811> A_IWL<12810> A_IWL<12809> A_IWL<12808> A_IWL<12807> A_IWL<12806> A_IWL<12805> A_IWL<12804> A_IWL<12803> A_IWL<12802> A_IWL<12801> A_IWL<12800> A_IWL<13311> A_IWL<13310> A_IWL<13309> A_IWL<13308> A_IWL<13307> A_IWL<13306> A_IWL<13305> A_IWL<13304> A_IWL<13303> A_IWL<13302> A_IWL<13301> A_IWL<13300> A_IWL<13299> A_IWL<13298> A_IWL<13297> A_IWL<13296> A_IWL<13295> A_IWL<13294> A_IWL<13293> A_IWL<13292> A_IWL<13291> A_IWL<13290> A_IWL<13289> A_IWL<13288> A_IWL<13287> A_IWL<13286> A_IWL<13285> A_IWL<13284> A_IWL<13283> A_IWL<13282> A_IWL<13281> A_IWL<13280> A_IWL<13279> A_IWL<13278> A_IWL<13277> A_IWL<13276> A_IWL<13275> A_IWL<13274> A_IWL<13273> A_IWL<13272> A_IWL<13271> A_IWL<13270> A_IWL<13269> A_IWL<13268> A_IWL<13267> A_IWL<13266> A_IWL<13265> A_IWL<13264> A_IWL<13263> A_IWL<13262> A_IWL<13261> A_IWL<13260> A_IWL<13259> A_IWL<13258> A_IWL<13257> A_IWL<13256> A_IWL<13255> A_IWL<13254> A_IWL<13253> A_IWL<13252> A_IWL<13251> A_IWL<13250> A_IWL<13249> A_IWL<13248> A_IWL<13247> A_IWL<13246> A_IWL<13245> A_IWL<13244> A_IWL<13243> A_IWL<13242> A_IWL<13241> A_IWL<13240> A_IWL<13239> A_IWL<13238> A_IWL<13237> A_IWL<13236> A_IWL<13235> A_IWL<13234> A_IWL<13233> A_IWL<13232> A_IWL<13231> A_IWL<13230> A_IWL<13229> A_IWL<13228> A_IWL<13227> A_IWL<13226> A_IWL<13225> A_IWL<13224> A_IWL<13223> A_IWL<13222> A_IWL<13221> A_IWL<13220> A_IWL<13219> A_IWL<13218> A_IWL<13217> A_IWL<13216> A_IWL<13215> A_IWL<13214> A_IWL<13213> A_IWL<13212> A_IWL<13211> A_IWL<13210> A_IWL<13209> A_IWL<13208> A_IWL<13207> A_IWL<13206> A_IWL<13205> A_IWL<13204> A_IWL<13203> A_IWL<13202> A_IWL<13201> A_IWL<13200> A_IWL<13199> A_IWL<13198> A_IWL<13197> A_IWL<13196> A_IWL<13195> A_IWL<13194> A_IWL<13193> A_IWL<13192> A_IWL<13191> A_IWL<13190> A_IWL<13189> A_IWL<13188> A_IWL<13187> A_IWL<13186> A_IWL<13185> A_IWL<13184> A_IWL<13183> A_IWL<13182> A_IWL<13181> A_IWL<13180> A_IWL<13179> A_IWL<13178> A_IWL<13177> A_IWL<13176> A_IWL<13175> A_IWL<13174> A_IWL<13173> A_IWL<13172> A_IWL<13171> A_IWL<13170> A_IWL<13169> A_IWL<13168> A_IWL<13167> A_IWL<13166> A_IWL<13165> A_IWL<13164> A_IWL<13163> A_IWL<13162> A_IWL<13161> A_IWL<13160> A_IWL<13159> A_IWL<13158> A_IWL<13157> A_IWL<13156> A_IWL<13155> A_IWL<13154> A_IWL<13153> A_IWL<13152> A_IWL<13151> A_IWL<13150> A_IWL<13149> A_IWL<13148> A_IWL<13147> A_IWL<13146> A_IWL<13145> A_IWL<13144> A_IWL<13143> A_IWL<13142> A_IWL<13141> A_IWL<13140> A_IWL<13139> A_IWL<13138> A_IWL<13137> A_IWL<13136> A_IWL<13135> A_IWL<13134> A_IWL<13133> A_IWL<13132> A_IWL<13131> A_IWL<13130> A_IWL<13129> A_IWL<13128> A_IWL<13127> A_IWL<13126> A_IWL<13125> A_IWL<13124> A_IWL<13123> A_IWL<13122> A_IWL<13121> A_IWL<13120> A_IWL<13119> A_IWL<13118> A_IWL<13117> A_IWL<13116> A_IWL<13115> A_IWL<13114> A_IWL<13113> A_IWL<13112> A_IWL<13111> A_IWL<13110> A_IWL<13109> A_IWL<13108> A_IWL<13107> A_IWL<13106> A_IWL<13105> A_IWL<13104> A_IWL<13103> A_IWL<13102> A_IWL<13101> A_IWL<13100> A_IWL<13099> A_IWL<13098> A_IWL<13097> A_IWL<13096> A_IWL<13095> A_IWL<13094> A_IWL<13093> A_IWL<13092> A_IWL<13091> A_IWL<13090> A_IWL<13089> A_IWL<13088> A_IWL<13087> A_IWL<13086> A_IWL<13085> A_IWL<13084> A_IWL<13083> A_IWL<13082> A_IWL<13081> A_IWL<13080> A_IWL<13079> A_IWL<13078> A_IWL<13077> A_IWL<13076> A_IWL<13075> A_IWL<13074> A_IWL<13073> A_IWL<13072> A_IWL<13071> A_IWL<13070> A_IWL<13069> A_IWL<13068> A_IWL<13067> A_IWL<13066> A_IWL<13065> A_IWL<13064> A_IWL<13063> A_IWL<13062> A_IWL<13061> A_IWL<13060> A_IWL<13059> A_IWL<13058> A_IWL<13057> A_IWL<13056> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<50> A_BLC<101> A_BLC<100> A_BLC_TOP<101> A_BLC_TOP<100> A_BLT<101> A_BLT<100> A_BLT_TOP<101> A_BLT_TOP<100> A_IWL<12799> A_IWL<12798> A_IWL<12797> A_IWL<12796> A_IWL<12795> A_IWL<12794> A_IWL<12793> A_IWL<12792> A_IWL<12791> A_IWL<12790> A_IWL<12789> A_IWL<12788> A_IWL<12787> A_IWL<12786> A_IWL<12785> A_IWL<12784> A_IWL<12783> A_IWL<12782> A_IWL<12781> A_IWL<12780> A_IWL<12779> A_IWL<12778> A_IWL<12777> A_IWL<12776> A_IWL<12775> A_IWL<12774> A_IWL<12773> A_IWL<12772> A_IWL<12771> A_IWL<12770> A_IWL<12769> A_IWL<12768> A_IWL<12767> A_IWL<12766> A_IWL<12765> A_IWL<12764> A_IWL<12763> A_IWL<12762> A_IWL<12761> A_IWL<12760> A_IWL<12759> A_IWL<12758> A_IWL<12757> A_IWL<12756> A_IWL<12755> A_IWL<12754> A_IWL<12753> A_IWL<12752> A_IWL<12751> A_IWL<12750> A_IWL<12749> A_IWL<12748> A_IWL<12747> A_IWL<12746> A_IWL<12745> A_IWL<12744> A_IWL<12743> A_IWL<12742> A_IWL<12741> A_IWL<12740> A_IWL<12739> A_IWL<12738> A_IWL<12737> A_IWL<12736> A_IWL<12735> A_IWL<12734> A_IWL<12733> A_IWL<12732> A_IWL<12731> A_IWL<12730> A_IWL<12729> A_IWL<12728> A_IWL<12727> A_IWL<12726> A_IWL<12725> A_IWL<12724> A_IWL<12723> A_IWL<12722> A_IWL<12721> A_IWL<12720> A_IWL<12719> A_IWL<12718> A_IWL<12717> A_IWL<12716> A_IWL<12715> A_IWL<12714> A_IWL<12713> A_IWL<12712> A_IWL<12711> A_IWL<12710> A_IWL<12709> A_IWL<12708> A_IWL<12707> A_IWL<12706> A_IWL<12705> A_IWL<12704> A_IWL<12703> A_IWL<12702> A_IWL<12701> A_IWL<12700> A_IWL<12699> A_IWL<12698> A_IWL<12697> A_IWL<12696> A_IWL<12695> A_IWL<12694> A_IWL<12693> A_IWL<12692> A_IWL<12691> A_IWL<12690> A_IWL<12689> A_IWL<12688> A_IWL<12687> A_IWL<12686> A_IWL<12685> A_IWL<12684> A_IWL<12683> A_IWL<12682> A_IWL<12681> A_IWL<12680> A_IWL<12679> A_IWL<12678> A_IWL<12677> A_IWL<12676> A_IWL<12675> A_IWL<12674> A_IWL<12673> A_IWL<12672> A_IWL<12671> A_IWL<12670> A_IWL<12669> A_IWL<12668> A_IWL<12667> A_IWL<12666> A_IWL<12665> A_IWL<12664> A_IWL<12663> A_IWL<12662> A_IWL<12661> A_IWL<12660> A_IWL<12659> A_IWL<12658> A_IWL<12657> A_IWL<12656> A_IWL<12655> A_IWL<12654> A_IWL<12653> A_IWL<12652> A_IWL<12651> A_IWL<12650> A_IWL<12649> A_IWL<12648> A_IWL<12647> A_IWL<12646> A_IWL<12645> A_IWL<12644> A_IWL<12643> A_IWL<12642> A_IWL<12641> A_IWL<12640> A_IWL<12639> A_IWL<12638> A_IWL<12637> A_IWL<12636> A_IWL<12635> A_IWL<12634> A_IWL<12633> A_IWL<12632> A_IWL<12631> A_IWL<12630> A_IWL<12629> A_IWL<12628> A_IWL<12627> A_IWL<12626> A_IWL<12625> A_IWL<12624> A_IWL<12623> A_IWL<12622> A_IWL<12621> A_IWL<12620> A_IWL<12619> A_IWL<12618> A_IWL<12617> A_IWL<12616> A_IWL<12615> A_IWL<12614> A_IWL<12613> A_IWL<12612> A_IWL<12611> A_IWL<12610> A_IWL<12609> A_IWL<12608> A_IWL<12607> A_IWL<12606> A_IWL<12605> A_IWL<12604> A_IWL<12603> A_IWL<12602> A_IWL<12601> A_IWL<12600> A_IWL<12599> A_IWL<12598> A_IWL<12597> A_IWL<12596> A_IWL<12595> A_IWL<12594> A_IWL<12593> A_IWL<12592> A_IWL<12591> A_IWL<12590> A_IWL<12589> A_IWL<12588> A_IWL<12587> A_IWL<12586> A_IWL<12585> A_IWL<12584> A_IWL<12583> A_IWL<12582> A_IWL<12581> A_IWL<12580> A_IWL<12579> A_IWL<12578> A_IWL<12577> A_IWL<12576> A_IWL<12575> A_IWL<12574> A_IWL<12573> A_IWL<12572> A_IWL<12571> A_IWL<12570> A_IWL<12569> A_IWL<12568> A_IWL<12567> A_IWL<12566> A_IWL<12565> A_IWL<12564> A_IWL<12563> A_IWL<12562> A_IWL<12561> A_IWL<12560> A_IWL<12559> A_IWL<12558> A_IWL<12557> A_IWL<12556> A_IWL<12555> A_IWL<12554> A_IWL<12553> A_IWL<12552> A_IWL<12551> A_IWL<12550> A_IWL<12549> A_IWL<12548> A_IWL<12547> A_IWL<12546> A_IWL<12545> A_IWL<12544> A_IWL<13055> A_IWL<13054> A_IWL<13053> A_IWL<13052> A_IWL<13051> A_IWL<13050> A_IWL<13049> A_IWL<13048> A_IWL<13047> A_IWL<13046> A_IWL<13045> A_IWL<13044> A_IWL<13043> A_IWL<13042> A_IWL<13041> A_IWL<13040> A_IWL<13039> A_IWL<13038> A_IWL<13037> A_IWL<13036> A_IWL<13035> A_IWL<13034> A_IWL<13033> A_IWL<13032> A_IWL<13031> A_IWL<13030> A_IWL<13029> A_IWL<13028> A_IWL<13027> A_IWL<13026> A_IWL<13025> A_IWL<13024> A_IWL<13023> A_IWL<13022> A_IWL<13021> A_IWL<13020> A_IWL<13019> A_IWL<13018> A_IWL<13017> A_IWL<13016> A_IWL<13015> A_IWL<13014> A_IWL<13013> A_IWL<13012> A_IWL<13011> A_IWL<13010> A_IWL<13009> A_IWL<13008> A_IWL<13007> A_IWL<13006> A_IWL<13005> A_IWL<13004> A_IWL<13003> A_IWL<13002> A_IWL<13001> A_IWL<13000> A_IWL<12999> A_IWL<12998> A_IWL<12997> A_IWL<12996> A_IWL<12995> A_IWL<12994> A_IWL<12993> A_IWL<12992> A_IWL<12991> A_IWL<12990> A_IWL<12989> A_IWL<12988> A_IWL<12987> A_IWL<12986> A_IWL<12985> A_IWL<12984> A_IWL<12983> A_IWL<12982> A_IWL<12981> A_IWL<12980> A_IWL<12979> A_IWL<12978> A_IWL<12977> A_IWL<12976> A_IWL<12975> A_IWL<12974> A_IWL<12973> A_IWL<12972> A_IWL<12971> A_IWL<12970> A_IWL<12969> A_IWL<12968> A_IWL<12967> A_IWL<12966> A_IWL<12965> A_IWL<12964> A_IWL<12963> A_IWL<12962> A_IWL<12961> A_IWL<12960> A_IWL<12959> A_IWL<12958> A_IWL<12957> A_IWL<12956> A_IWL<12955> A_IWL<12954> A_IWL<12953> A_IWL<12952> A_IWL<12951> A_IWL<12950> A_IWL<12949> A_IWL<12948> A_IWL<12947> A_IWL<12946> A_IWL<12945> A_IWL<12944> A_IWL<12943> A_IWL<12942> A_IWL<12941> A_IWL<12940> A_IWL<12939> A_IWL<12938> A_IWL<12937> A_IWL<12936> A_IWL<12935> A_IWL<12934> A_IWL<12933> A_IWL<12932> A_IWL<12931> A_IWL<12930> A_IWL<12929> A_IWL<12928> A_IWL<12927> A_IWL<12926> A_IWL<12925> A_IWL<12924> A_IWL<12923> A_IWL<12922> A_IWL<12921> A_IWL<12920> A_IWL<12919> A_IWL<12918> A_IWL<12917> A_IWL<12916> A_IWL<12915> A_IWL<12914> A_IWL<12913> A_IWL<12912> A_IWL<12911> A_IWL<12910> A_IWL<12909> A_IWL<12908> A_IWL<12907> A_IWL<12906> A_IWL<12905> A_IWL<12904> A_IWL<12903> A_IWL<12902> A_IWL<12901> A_IWL<12900> A_IWL<12899> A_IWL<12898> A_IWL<12897> A_IWL<12896> A_IWL<12895> A_IWL<12894> A_IWL<12893> A_IWL<12892> A_IWL<12891> A_IWL<12890> A_IWL<12889> A_IWL<12888> A_IWL<12887> A_IWL<12886> A_IWL<12885> A_IWL<12884> A_IWL<12883> A_IWL<12882> A_IWL<12881> A_IWL<12880> A_IWL<12879> A_IWL<12878> A_IWL<12877> A_IWL<12876> A_IWL<12875> A_IWL<12874> A_IWL<12873> A_IWL<12872> A_IWL<12871> A_IWL<12870> A_IWL<12869> A_IWL<12868> A_IWL<12867> A_IWL<12866> A_IWL<12865> A_IWL<12864> A_IWL<12863> A_IWL<12862> A_IWL<12861> A_IWL<12860> A_IWL<12859> A_IWL<12858> A_IWL<12857> A_IWL<12856> A_IWL<12855> A_IWL<12854> A_IWL<12853> A_IWL<12852> A_IWL<12851> A_IWL<12850> A_IWL<12849> A_IWL<12848> A_IWL<12847> A_IWL<12846> A_IWL<12845> A_IWL<12844> A_IWL<12843> A_IWL<12842> A_IWL<12841> A_IWL<12840> A_IWL<12839> A_IWL<12838> A_IWL<12837> A_IWL<12836> A_IWL<12835> A_IWL<12834> A_IWL<12833> A_IWL<12832> A_IWL<12831> A_IWL<12830> A_IWL<12829> A_IWL<12828> A_IWL<12827> A_IWL<12826> A_IWL<12825> A_IWL<12824> A_IWL<12823> A_IWL<12822> A_IWL<12821> A_IWL<12820> A_IWL<12819> A_IWL<12818> A_IWL<12817> A_IWL<12816> A_IWL<12815> A_IWL<12814> A_IWL<12813> A_IWL<12812> A_IWL<12811> A_IWL<12810> A_IWL<12809> A_IWL<12808> A_IWL<12807> A_IWL<12806> A_IWL<12805> A_IWL<12804> A_IWL<12803> A_IWL<12802> A_IWL<12801> A_IWL<12800> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<49> A_BLC<99> A_BLC<98> A_BLC_TOP<99> A_BLC_TOP<98> A_BLT<99> A_BLT<98> A_BLT_TOP<99> A_BLT_TOP<98> A_IWL<12543> A_IWL<12542> A_IWL<12541> A_IWL<12540> A_IWL<12539> A_IWL<12538> A_IWL<12537> A_IWL<12536> A_IWL<12535> A_IWL<12534> A_IWL<12533> A_IWL<12532> A_IWL<12531> A_IWL<12530> A_IWL<12529> A_IWL<12528> A_IWL<12527> A_IWL<12526> A_IWL<12525> A_IWL<12524> A_IWL<12523> A_IWL<12522> A_IWL<12521> A_IWL<12520> A_IWL<12519> A_IWL<12518> A_IWL<12517> A_IWL<12516> A_IWL<12515> A_IWL<12514> A_IWL<12513> A_IWL<12512> A_IWL<12511> A_IWL<12510> A_IWL<12509> A_IWL<12508> A_IWL<12507> A_IWL<12506> A_IWL<12505> A_IWL<12504> A_IWL<12503> A_IWL<12502> A_IWL<12501> A_IWL<12500> A_IWL<12499> A_IWL<12498> A_IWL<12497> A_IWL<12496> A_IWL<12495> A_IWL<12494> A_IWL<12493> A_IWL<12492> A_IWL<12491> A_IWL<12490> A_IWL<12489> A_IWL<12488> A_IWL<12487> A_IWL<12486> A_IWL<12485> A_IWL<12484> A_IWL<12483> A_IWL<12482> A_IWL<12481> A_IWL<12480> A_IWL<12479> A_IWL<12478> A_IWL<12477> A_IWL<12476> A_IWL<12475> A_IWL<12474> A_IWL<12473> A_IWL<12472> A_IWL<12471> A_IWL<12470> A_IWL<12469> A_IWL<12468> A_IWL<12467> A_IWL<12466> A_IWL<12465> A_IWL<12464> A_IWL<12463> A_IWL<12462> A_IWL<12461> A_IWL<12460> A_IWL<12459> A_IWL<12458> A_IWL<12457> A_IWL<12456> A_IWL<12455> A_IWL<12454> A_IWL<12453> A_IWL<12452> A_IWL<12451> A_IWL<12450> A_IWL<12449> A_IWL<12448> A_IWL<12447> A_IWL<12446> A_IWL<12445> A_IWL<12444> A_IWL<12443> A_IWL<12442> A_IWL<12441> A_IWL<12440> A_IWL<12439> A_IWL<12438> A_IWL<12437> A_IWL<12436> A_IWL<12435> A_IWL<12434> A_IWL<12433> A_IWL<12432> A_IWL<12431> A_IWL<12430> A_IWL<12429> A_IWL<12428> A_IWL<12427> A_IWL<12426> A_IWL<12425> A_IWL<12424> A_IWL<12423> A_IWL<12422> A_IWL<12421> A_IWL<12420> A_IWL<12419> A_IWL<12418> A_IWL<12417> A_IWL<12416> A_IWL<12415> A_IWL<12414> A_IWL<12413> A_IWL<12412> A_IWL<12411> A_IWL<12410> A_IWL<12409> A_IWL<12408> A_IWL<12407> A_IWL<12406> A_IWL<12405> A_IWL<12404> A_IWL<12403> A_IWL<12402> A_IWL<12401> A_IWL<12400> A_IWL<12399> A_IWL<12398> A_IWL<12397> A_IWL<12396> A_IWL<12395> A_IWL<12394> A_IWL<12393> A_IWL<12392> A_IWL<12391> A_IWL<12390> A_IWL<12389> A_IWL<12388> A_IWL<12387> A_IWL<12386> A_IWL<12385> A_IWL<12384> A_IWL<12383> A_IWL<12382> A_IWL<12381> A_IWL<12380> A_IWL<12379> A_IWL<12378> A_IWL<12377> A_IWL<12376> A_IWL<12375> A_IWL<12374> A_IWL<12373> A_IWL<12372> A_IWL<12371> A_IWL<12370> A_IWL<12369> A_IWL<12368> A_IWL<12367> A_IWL<12366> A_IWL<12365> A_IWL<12364> A_IWL<12363> A_IWL<12362> A_IWL<12361> A_IWL<12360> A_IWL<12359> A_IWL<12358> A_IWL<12357> A_IWL<12356> A_IWL<12355> A_IWL<12354> A_IWL<12353> A_IWL<12352> A_IWL<12351> A_IWL<12350> A_IWL<12349> A_IWL<12348> A_IWL<12347> A_IWL<12346> A_IWL<12345> A_IWL<12344> A_IWL<12343> A_IWL<12342> A_IWL<12341> A_IWL<12340> A_IWL<12339> A_IWL<12338> A_IWL<12337> A_IWL<12336> A_IWL<12335> A_IWL<12334> A_IWL<12333> A_IWL<12332> A_IWL<12331> A_IWL<12330> A_IWL<12329> A_IWL<12328> A_IWL<12327> A_IWL<12326> A_IWL<12325> A_IWL<12324> A_IWL<12323> A_IWL<12322> A_IWL<12321> A_IWL<12320> A_IWL<12319> A_IWL<12318> A_IWL<12317> A_IWL<12316> A_IWL<12315> A_IWL<12314> A_IWL<12313> A_IWL<12312> A_IWL<12311> A_IWL<12310> A_IWL<12309> A_IWL<12308> A_IWL<12307> A_IWL<12306> A_IWL<12305> A_IWL<12304> A_IWL<12303> A_IWL<12302> A_IWL<12301> A_IWL<12300> A_IWL<12299> A_IWL<12298> A_IWL<12297> A_IWL<12296> A_IWL<12295> A_IWL<12294> A_IWL<12293> A_IWL<12292> A_IWL<12291> A_IWL<12290> A_IWL<12289> A_IWL<12288> A_IWL<12799> A_IWL<12798> A_IWL<12797> A_IWL<12796> A_IWL<12795> A_IWL<12794> A_IWL<12793> A_IWL<12792> A_IWL<12791> A_IWL<12790> A_IWL<12789> A_IWL<12788> A_IWL<12787> A_IWL<12786> A_IWL<12785> A_IWL<12784> A_IWL<12783> A_IWL<12782> A_IWL<12781> A_IWL<12780> A_IWL<12779> A_IWL<12778> A_IWL<12777> A_IWL<12776> A_IWL<12775> A_IWL<12774> A_IWL<12773> A_IWL<12772> A_IWL<12771> A_IWL<12770> A_IWL<12769> A_IWL<12768> A_IWL<12767> A_IWL<12766> A_IWL<12765> A_IWL<12764> A_IWL<12763> A_IWL<12762> A_IWL<12761> A_IWL<12760> A_IWL<12759> A_IWL<12758> A_IWL<12757> A_IWL<12756> A_IWL<12755> A_IWL<12754> A_IWL<12753> A_IWL<12752> A_IWL<12751> A_IWL<12750> A_IWL<12749> A_IWL<12748> A_IWL<12747> A_IWL<12746> A_IWL<12745> A_IWL<12744> A_IWL<12743> A_IWL<12742> A_IWL<12741> A_IWL<12740> A_IWL<12739> A_IWL<12738> A_IWL<12737> A_IWL<12736> A_IWL<12735> A_IWL<12734> A_IWL<12733> A_IWL<12732> A_IWL<12731> A_IWL<12730> A_IWL<12729> A_IWL<12728> A_IWL<12727> A_IWL<12726> A_IWL<12725> A_IWL<12724> A_IWL<12723> A_IWL<12722> A_IWL<12721> A_IWL<12720> A_IWL<12719> A_IWL<12718> A_IWL<12717> A_IWL<12716> A_IWL<12715> A_IWL<12714> A_IWL<12713> A_IWL<12712> A_IWL<12711> A_IWL<12710> A_IWL<12709> A_IWL<12708> A_IWL<12707> A_IWL<12706> A_IWL<12705> A_IWL<12704> A_IWL<12703> A_IWL<12702> A_IWL<12701> A_IWL<12700> A_IWL<12699> A_IWL<12698> A_IWL<12697> A_IWL<12696> A_IWL<12695> A_IWL<12694> A_IWL<12693> A_IWL<12692> A_IWL<12691> A_IWL<12690> A_IWL<12689> A_IWL<12688> A_IWL<12687> A_IWL<12686> A_IWL<12685> A_IWL<12684> A_IWL<12683> A_IWL<12682> A_IWL<12681> A_IWL<12680> A_IWL<12679> A_IWL<12678> A_IWL<12677> A_IWL<12676> A_IWL<12675> A_IWL<12674> A_IWL<12673> A_IWL<12672> A_IWL<12671> A_IWL<12670> A_IWL<12669> A_IWL<12668> A_IWL<12667> A_IWL<12666> A_IWL<12665> A_IWL<12664> A_IWL<12663> A_IWL<12662> A_IWL<12661> A_IWL<12660> A_IWL<12659> A_IWL<12658> A_IWL<12657> A_IWL<12656> A_IWL<12655> A_IWL<12654> A_IWL<12653> A_IWL<12652> A_IWL<12651> A_IWL<12650> A_IWL<12649> A_IWL<12648> A_IWL<12647> A_IWL<12646> A_IWL<12645> A_IWL<12644> A_IWL<12643> A_IWL<12642> A_IWL<12641> A_IWL<12640> A_IWL<12639> A_IWL<12638> A_IWL<12637> A_IWL<12636> A_IWL<12635> A_IWL<12634> A_IWL<12633> A_IWL<12632> A_IWL<12631> A_IWL<12630> A_IWL<12629> A_IWL<12628> A_IWL<12627> A_IWL<12626> A_IWL<12625> A_IWL<12624> A_IWL<12623> A_IWL<12622> A_IWL<12621> A_IWL<12620> A_IWL<12619> A_IWL<12618> A_IWL<12617> A_IWL<12616> A_IWL<12615> A_IWL<12614> A_IWL<12613> A_IWL<12612> A_IWL<12611> A_IWL<12610> A_IWL<12609> A_IWL<12608> A_IWL<12607> A_IWL<12606> A_IWL<12605> A_IWL<12604> A_IWL<12603> A_IWL<12602> A_IWL<12601> A_IWL<12600> A_IWL<12599> A_IWL<12598> A_IWL<12597> A_IWL<12596> A_IWL<12595> A_IWL<12594> A_IWL<12593> A_IWL<12592> A_IWL<12591> A_IWL<12590> A_IWL<12589> A_IWL<12588> A_IWL<12587> A_IWL<12586> A_IWL<12585> A_IWL<12584> A_IWL<12583> A_IWL<12582> A_IWL<12581> A_IWL<12580> A_IWL<12579> A_IWL<12578> A_IWL<12577> A_IWL<12576> A_IWL<12575> A_IWL<12574> A_IWL<12573> A_IWL<12572> A_IWL<12571> A_IWL<12570> A_IWL<12569> A_IWL<12568> A_IWL<12567> A_IWL<12566> A_IWL<12565> A_IWL<12564> A_IWL<12563> A_IWL<12562> A_IWL<12561> A_IWL<12560> A_IWL<12559> A_IWL<12558> A_IWL<12557> A_IWL<12556> A_IWL<12555> A_IWL<12554> A_IWL<12553> A_IWL<12552> A_IWL<12551> A_IWL<12550> A_IWL<12549> A_IWL<12548> A_IWL<12547> A_IWL<12546> A_IWL<12545> A_IWL<12544> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<48> A_BLC<97> A_BLC<96> A_BLC_TOP<97> A_BLC_TOP<96> A_BLT<97> A_BLT<96> A_BLT_TOP<97> A_BLT_TOP<96> A_IWL<12287> A_IWL<12286> A_IWL<12285> A_IWL<12284> A_IWL<12283> A_IWL<12282> A_IWL<12281> A_IWL<12280> A_IWL<12279> A_IWL<12278> A_IWL<12277> A_IWL<12276> A_IWL<12275> A_IWL<12274> A_IWL<12273> A_IWL<12272> A_IWL<12271> A_IWL<12270> A_IWL<12269> A_IWL<12268> A_IWL<12267> A_IWL<12266> A_IWL<12265> A_IWL<12264> A_IWL<12263> A_IWL<12262> A_IWL<12261> A_IWL<12260> A_IWL<12259> A_IWL<12258> A_IWL<12257> A_IWL<12256> A_IWL<12255> A_IWL<12254> A_IWL<12253> A_IWL<12252> A_IWL<12251> A_IWL<12250> A_IWL<12249> A_IWL<12248> A_IWL<12247> A_IWL<12246> A_IWL<12245> A_IWL<12244> A_IWL<12243> A_IWL<12242> A_IWL<12241> A_IWL<12240> A_IWL<12239> A_IWL<12238> A_IWL<12237> A_IWL<12236> A_IWL<12235> A_IWL<12234> A_IWL<12233> A_IWL<12232> A_IWL<12231> A_IWL<12230> A_IWL<12229> A_IWL<12228> A_IWL<12227> A_IWL<12226> A_IWL<12225> A_IWL<12224> A_IWL<12223> A_IWL<12222> A_IWL<12221> A_IWL<12220> A_IWL<12219> A_IWL<12218> A_IWL<12217> A_IWL<12216> A_IWL<12215> A_IWL<12214> A_IWL<12213> A_IWL<12212> A_IWL<12211> A_IWL<12210> A_IWL<12209> A_IWL<12208> A_IWL<12207> A_IWL<12206> A_IWL<12205> A_IWL<12204> A_IWL<12203> A_IWL<12202> A_IWL<12201> A_IWL<12200> A_IWL<12199> A_IWL<12198> A_IWL<12197> A_IWL<12196> A_IWL<12195> A_IWL<12194> A_IWL<12193> A_IWL<12192> A_IWL<12191> A_IWL<12190> A_IWL<12189> A_IWL<12188> A_IWL<12187> A_IWL<12186> A_IWL<12185> A_IWL<12184> A_IWL<12183> A_IWL<12182> A_IWL<12181> A_IWL<12180> A_IWL<12179> A_IWL<12178> A_IWL<12177> A_IWL<12176> A_IWL<12175> A_IWL<12174> A_IWL<12173> A_IWL<12172> A_IWL<12171> A_IWL<12170> A_IWL<12169> A_IWL<12168> A_IWL<12167> A_IWL<12166> A_IWL<12165> A_IWL<12164> A_IWL<12163> A_IWL<12162> A_IWL<12161> A_IWL<12160> A_IWL<12159> A_IWL<12158> A_IWL<12157> A_IWL<12156> A_IWL<12155> A_IWL<12154> A_IWL<12153> A_IWL<12152> A_IWL<12151> A_IWL<12150> A_IWL<12149> A_IWL<12148> A_IWL<12147> A_IWL<12146> A_IWL<12145> A_IWL<12144> A_IWL<12143> A_IWL<12142> A_IWL<12141> A_IWL<12140> A_IWL<12139> A_IWL<12138> A_IWL<12137> A_IWL<12136> A_IWL<12135> A_IWL<12134> A_IWL<12133> A_IWL<12132> A_IWL<12131> A_IWL<12130> A_IWL<12129> A_IWL<12128> A_IWL<12127> A_IWL<12126> A_IWL<12125> A_IWL<12124> A_IWL<12123> A_IWL<12122> A_IWL<12121> A_IWL<12120> A_IWL<12119> A_IWL<12118> A_IWL<12117> A_IWL<12116> A_IWL<12115> A_IWL<12114> A_IWL<12113> A_IWL<12112> A_IWL<12111> A_IWL<12110> A_IWL<12109> A_IWL<12108> A_IWL<12107> A_IWL<12106> A_IWL<12105> A_IWL<12104> A_IWL<12103> A_IWL<12102> A_IWL<12101> A_IWL<12100> A_IWL<12099> A_IWL<12098> A_IWL<12097> A_IWL<12096> A_IWL<12095> A_IWL<12094> A_IWL<12093> A_IWL<12092> A_IWL<12091> A_IWL<12090> A_IWL<12089> A_IWL<12088> A_IWL<12087> A_IWL<12086> A_IWL<12085> A_IWL<12084> A_IWL<12083> A_IWL<12082> A_IWL<12081> A_IWL<12080> A_IWL<12079> A_IWL<12078> A_IWL<12077> A_IWL<12076> A_IWL<12075> A_IWL<12074> A_IWL<12073> A_IWL<12072> A_IWL<12071> A_IWL<12070> A_IWL<12069> A_IWL<12068> A_IWL<12067> A_IWL<12066> A_IWL<12065> A_IWL<12064> A_IWL<12063> A_IWL<12062> A_IWL<12061> A_IWL<12060> A_IWL<12059> A_IWL<12058> A_IWL<12057> A_IWL<12056> A_IWL<12055> A_IWL<12054> A_IWL<12053> A_IWL<12052> A_IWL<12051> A_IWL<12050> A_IWL<12049> A_IWL<12048> A_IWL<12047> A_IWL<12046> A_IWL<12045> A_IWL<12044> A_IWL<12043> A_IWL<12042> A_IWL<12041> A_IWL<12040> A_IWL<12039> A_IWL<12038> A_IWL<12037> A_IWL<12036> A_IWL<12035> A_IWL<12034> A_IWL<12033> A_IWL<12032> A_IWL<12543> A_IWL<12542> A_IWL<12541> A_IWL<12540> A_IWL<12539> A_IWL<12538> A_IWL<12537> A_IWL<12536> A_IWL<12535> A_IWL<12534> A_IWL<12533> A_IWL<12532> A_IWL<12531> A_IWL<12530> A_IWL<12529> A_IWL<12528> A_IWL<12527> A_IWL<12526> A_IWL<12525> A_IWL<12524> A_IWL<12523> A_IWL<12522> A_IWL<12521> A_IWL<12520> A_IWL<12519> A_IWL<12518> A_IWL<12517> A_IWL<12516> A_IWL<12515> A_IWL<12514> A_IWL<12513> A_IWL<12512> A_IWL<12511> A_IWL<12510> A_IWL<12509> A_IWL<12508> A_IWL<12507> A_IWL<12506> A_IWL<12505> A_IWL<12504> A_IWL<12503> A_IWL<12502> A_IWL<12501> A_IWL<12500> A_IWL<12499> A_IWL<12498> A_IWL<12497> A_IWL<12496> A_IWL<12495> A_IWL<12494> A_IWL<12493> A_IWL<12492> A_IWL<12491> A_IWL<12490> A_IWL<12489> A_IWL<12488> A_IWL<12487> A_IWL<12486> A_IWL<12485> A_IWL<12484> A_IWL<12483> A_IWL<12482> A_IWL<12481> A_IWL<12480> A_IWL<12479> A_IWL<12478> A_IWL<12477> A_IWL<12476> A_IWL<12475> A_IWL<12474> A_IWL<12473> A_IWL<12472> A_IWL<12471> A_IWL<12470> A_IWL<12469> A_IWL<12468> A_IWL<12467> A_IWL<12466> A_IWL<12465> A_IWL<12464> A_IWL<12463> A_IWL<12462> A_IWL<12461> A_IWL<12460> A_IWL<12459> A_IWL<12458> A_IWL<12457> A_IWL<12456> A_IWL<12455> A_IWL<12454> A_IWL<12453> A_IWL<12452> A_IWL<12451> A_IWL<12450> A_IWL<12449> A_IWL<12448> A_IWL<12447> A_IWL<12446> A_IWL<12445> A_IWL<12444> A_IWL<12443> A_IWL<12442> A_IWL<12441> A_IWL<12440> A_IWL<12439> A_IWL<12438> A_IWL<12437> A_IWL<12436> A_IWL<12435> A_IWL<12434> A_IWL<12433> A_IWL<12432> A_IWL<12431> A_IWL<12430> A_IWL<12429> A_IWL<12428> A_IWL<12427> A_IWL<12426> A_IWL<12425> A_IWL<12424> A_IWL<12423> A_IWL<12422> A_IWL<12421> A_IWL<12420> A_IWL<12419> A_IWL<12418> A_IWL<12417> A_IWL<12416> A_IWL<12415> A_IWL<12414> A_IWL<12413> A_IWL<12412> A_IWL<12411> A_IWL<12410> A_IWL<12409> A_IWL<12408> A_IWL<12407> A_IWL<12406> A_IWL<12405> A_IWL<12404> A_IWL<12403> A_IWL<12402> A_IWL<12401> A_IWL<12400> A_IWL<12399> A_IWL<12398> A_IWL<12397> A_IWL<12396> A_IWL<12395> A_IWL<12394> A_IWL<12393> A_IWL<12392> A_IWL<12391> A_IWL<12390> A_IWL<12389> A_IWL<12388> A_IWL<12387> A_IWL<12386> A_IWL<12385> A_IWL<12384> A_IWL<12383> A_IWL<12382> A_IWL<12381> A_IWL<12380> A_IWL<12379> A_IWL<12378> A_IWL<12377> A_IWL<12376> A_IWL<12375> A_IWL<12374> A_IWL<12373> A_IWL<12372> A_IWL<12371> A_IWL<12370> A_IWL<12369> A_IWL<12368> A_IWL<12367> A_IWL<12366> A_IWL<12365> A_IWL<12364> A_IWL<12363> A_IWL<12362> A_IWL<12361> A_IWL<12360> A_IWL<12359> A_IWL<12358> A_IWL<12357> A_IWL<12356> A_IWL<12355> A_IWL<12354> A_IWL<12353> A_IWL<12352> A_IWL<12351> A_IWL<12350> A_IWL<12349> A_IWL<12348> A_IWL<12347> A_IWL<12346> A_IWL<12345> A_IWL<12344> A_IWL<12343> A_IWL<12342> A_IWL<12341> A_IWL<12340> A_IWL<12339> A_IWL<12338> A_IWL<12337> A_IWL<12336> A_IWL<12335> A_IWL<12334> A_IWL<12333> A_IWL<12332> A_IWL<12331> A_IWL<12330> A_IWL<12329> A_IWL<12328> A_IWL<12327> A_IWL<12326> A_IWL<12325> A_IWL<12324> A_IWL<12323> A_IWL<12322> A_IWL<12321> A_IWL<12320> A_IWL<12319> A_IWL<12318> A_IWL<12317> A_IWL<12316> A_IWL<12315> A_IWL<12314> A_IWL<12313> A_IWL<12312> A_IWL<12311> A_IWL<12310> A_IWL<12309> A_IWL<12308> A_IWL<12307> A_IWL<12306> A_IWL<12305> A_IWL<12304> A_IWL<12303> A_IWL<12302> A_IWL<12301> A_IWL<12300> A_IWL<12299> A_IWL<12298> A_IWL<12297> A_IWL<12296> A_IWL<12295> A_IWL<12294> A_IWL<12293> A_IWL<12292> A_IWL<12291> A_IWL<12290> A_IWL<12289> A_IWL<12288> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<47> A_BLC<95> A_BLC<94> A_BLC_TOP<95> A_BLC_TOP<94> A_BLT<95> A_BLT<94> A_BLT_TOP<95> A_BLT_TOP<94> A_IWL<12031> A_IWL<12030> A_IWL<12029> A_IWL<12028> A_IWL<12027> A_IWL<12026> A_IWL<12025> A_IWL<12024> A_IWL<12023> A_IWL<12022> A_IWL<12021> A_IWL<12020> A_IWL<12019> A_IWL<12018> A_IWL<12017> A_IWL<12016> A_IWL<12015> A_IWL<12014> A_IWL<12013> A_IWL<12012> A_IWL<12011> A_IWL<12010> A_IWL<12009> A_IWL<12008> A_IWL<12007> A_IWL<12006> A_IWL<12005> A_IWL<12004> A_IWL<12003> A_IWL<12002> A_IWL<12001> A_IWL<12000> A_IWL<11999> A_IWL<11998> A_IWL<11997> A_IWL<11996> A_IWL<11995> A_IWL<11994> A_IWL<11993> A_IWL<11992> A_IWL<11991> A_IWL<11990> A_IWL<11989> A_IWL<11988> A_IWL<11987> A_IWL<11986> A_IWL<11985> A_IWL<11984> A_IWL<11983> A_IWL<11982> A_IWL<11981> A_IWL<11980> A_IWL<11979> A_IWL<11978> A_IWL<11977> A_IWL<11976> A_IWL<11975> A_IWL<11974> A_IWL<11973> A_IWL<11972> A_IWL<11971> A_IWL<11970> A_IWL<11969> A_IWL<11968> A_IWL<11967> A_IWL<11966> A_IWL<11965> A_IWL<11964> A_IWL<11963> A_IWL<11962> A_IWL<11961> A_IWL<11960> A_IWL<11959> A_IWL<11958> A_IWL<11957> A_IWL<11956> A_IWL<11955> A_IWL<11954> A_IWL<11953> A_IWL<11952> A_IWL<11951> A_IWL<11950> A_IWL<11949> A_IWL<11948> A_IWL<11947> A_IWL<11946> A_IWL<11945> A_IWL<11944> A_IWL<11943> A_IWL<11942> A_IWL<11941> A_IWL<11940> A_IWL<11939> A_IWL<11938> A_IWL<11937> A_IWL<11936> A_IWL<11935> A_IWL<11934> A_IWL<11933> A_IWL<11932> A_IWL<11931> A_IWL<11930> A_IWL<11929> A_IWL<11928> A_IWL<11927> A_IWL<11926> A_IWL<11925> A_IWL<11924> A_IWL<11923> A_IWL<11922> A_IWL<11921> A_IWL<11920> A_IWL<11919> A_IWL<11918> A_IWL<11917> A_IWL<11916> A_IWL<11915> A_IWL<11914> A_IWL<11913> A_IWL<11912> A_IWL<11911> A_IWL<11910> A_IWL<11909> A_IWL<11908> A_IWL<11907> A_IWL<11906> A_IWL<11905> A_IWL<11904> A_IWL<11903> A_IWL<11902> A_IWL<11901> A_IWL<11900> A_IWL<11899> A_IWL<11898> A_IWL<11897> A_IWL<11896> A_IWL<11895> A_IWL<11894> A_IWL<11893> A_IWL<11892> A_IWL<11891> A_IWL<11890> A_IWL<11889> A_IWL<11888> A_IWL<11887> A_IWL<11886> A_IWL<11885> A_IWL<11884> A_IWL<11883> A_IWL<11882> A_IWL<11881> A_IWL<11880> A_IWL<11879> A_IWL<11878> A_IWL<11877> A_IWL<11876> A_IWL<11875> A_IWL<11874> A_IWL<11873> A_IWL<11872> A_IWL<11871> A_IWL<11870> A_IWL<11869> A_IWL<11868> A_IWL<11867> A_IWL<11866> A_IWL<11865> A_IWL<11864> A_IWL<11863> A_IWL<11862> A_IWL<11861> A_IWL<11860> A_IWL<11859> A_IWL<11858> A_IWL<11857> A_IWL<11856> A_IWL<11855> A_IWL<11854> A_IWL<11853> A_IWL<11852> A_IWL<11851> A_IWL<11850> A_IWL<11849> A_IWL<11848> A_IWL<11847> A_IWL<11846> A_IWL<11845> A_IWL<11844> A_IWL<11843> A_IWL<11842> A_IWL<11841> A_IWL<11840> A_IWL<11839> A_IWL<11838> A_IWL<11837> A_IWL<11836> A_IWL<11835> A_IWL<11834> A_IWL<11833> A_IWL<11832> A_IWL<11831> A_IWL<11830> A_IWL<11829> A_IWL<11828> A_IWL<11827> A_IWL<11826> A_IWL<11825> A_IWL<11824> A_IWL<11823> A_IWL<11822> A_IWL<11821> A_IWL<11820> A_IWL<11819> A_IWL<11818> A_IWL<11817> A_IWL<11816> A_IWL<11815> A_IWL<11814> A_IWL<11813> A_IWL<11812> A_IWL<11811> A_IWL<11810> A_IWL<11809> A_IWL<11808> A_IWL<11807> A_IWL<11806> A_IWL<11805> A_IWL<11804> A_IWL<11803> A_IWL<11802> A_IWL<11801> A_IWL<11800> A_IWL<11799> A_IWL<11798> A_IWL<11797> A_IWL<11796> A_IWL<11795> A_IWL<11794> A_IWL<11793> A_IWL<11792> A_IWL<11791> A_IWL<11790> A_IWL<11789> A_IWL<11788> A_IWL<11787> A_IWL<11786> A_IWL<11785> A_IWL<11784> A_IWL<11783> A_IWL<11782> A_IWL<11781> A_IWL<11780> A_IWL<11779> A_IWL<11778> A_IWL<11777> A_IWL<11776> A_IWL<12287> A_IWL<12286> A_IWL<12285> A_IWL<12284> A_IWL<12283> A_IWL<12282> A_IWL<12281> A_IWL<12280> A_IWL<12279> A_IWL<12278> A_IWL<12277> A_IWL<12276> A_IWL<12275> A_IWL<12274> A_IWL<12273> A_IWL<12272> A_IWL<12271> A_IWL<12270> A_IWL<12269> A_IWL<12268> A_IWL<12267> A_IWL<12266> A_IWL<12265> A_IWL<12264> A_IWL<12263> A_IWL<12262> A_IWL<12261> A_IWL<12260> A_IWL<12259> A_IWL<12258> A_IWL<12257> A_IWL<12256> A_IWL<12255> A_IWL<12254> A_IWL<12253> A_IWL<12252> A_IWL<12251> A_IWL<12250> A_IWL<12249> A_IWL<12248> A_IWL<12247> A_IWL<12246> A_IWL<12245> A_IWL<12244> A_IWL<12243> A_IWL<12242> A_IWL<12241> A_IWL<12240> A_IWL<12239> A_IWL<12238> A_IWL<12237> A_IWL<12236> A_IWL<12235> A_IWL<12234> A_IWL<12233> A_IWL<12232> A_IWL<12231> A_IWL<12230> A_IWL<12229> A_IWL<12228> A_IWL<12227> A_IWL<12226> A_IWL<12225> A_IWL<12224> A_IWL<12223> A_IWL<12222> A_IWL<12221> A_IWL<12220> A_IWL<12219> A_IWL<12218> A_IWL<12217> A_IWL<12216> A_IWL<12215> A_IWL<12214> A_IWL<12213> A_IWL<12212> A_IWL<12211> A_IWL<12210> A_IWL<12209> A_IWL<12208> A_IWL<12207> A_IWL<12206> A_IWL<12205> A_IWL<12204> A_IWL<12203> A_IWL<12202> A_IWL<12201> A_IWL<12200> A_IWL<12199> A_IWL<12198> A_IWL<12197> A_IWL<12196> A_IWL<12195> A_IWL<12194> A_IWL<12193> A_IWL<12192> A_IWL<12191> A_IWL<12190> A_IWL<12189> A_IWL<12188> A_IWL<12187> A_IWL<12186> A_IWL<12185> A_IWL<12184> A_IWL<12183> A_IWL<12182> A_IWL<12181> A_IWL<12180> A_IWL<12179> A_IWL<12178> A_IWL<12177> A_IWL<12176> A_IWL<12175> A_IWL<12174> A_IWL<12173> A_IWL<12172> A_IWL<12171> A_IWL<12170> A_IWL<12169> A_IWL<12168> A_IWL<12167> A_IWL<12166> A_IWL<12165> A_IWL<12164> A_IWL<12163> A_IWL<12162> A_IWL<12161> A_IWL<12160> A_IWL<12159> A_IWL<12158> A_IWL<12157> A_IWL<12156> A_IWL<12155> A_IWL<12154> A_IWL<12153> A_IWL<12152> A_IWL<12151> A_IWL<12150> A_IWL<12149> A_IWL<12148> A_IWL<12147> A_IWL<12146> A_IWL<12145> A_IWL<12144> A_IWL<12143> A_IWL<12142> A_IWL<12141> A_IWL<12140> A_IWL<12139> A_IWL<12138> A_IWL<12137> A_IWL<12136> A_IWL<12135> A_IWL<12134> A_IWL<12133> A_IWL<12132> A_IWL<12131> A_IWL<12130> A_IWL<12129> A_IWL<12128> A_IWL<12127> A_IWL<12126> A_IWL<12125> A_IWL<12124> A_IWL<12123> A_IWL<12122> A_IWL<12121> A_IWL<12120> A_IWL<12119> A_IWL<12118> A_IWL<12117> A_IWL<12116> A_IWL<12115> A_IWL<12114> A_IWL<12113> A_IWL<12112> A_IWL<12111> A_IWL<12110> A_IWL<12109> A_IWL<12108> A_IWL<12107> A_IWL<12106> A_IWL<12105> A_IWL<12104> A_IWL<12103> A_IWL<12102> A_IWL<12101> A_IWL<12100> A_IWL<12099> A_IWL<12098> A_IWL<12097> A_IWL<12096> A_IWL<12095> A_IWL<12094> A_IWL<12093> A_IWL<12092> A_IWL<12091> A_IWL<12090> A_IWL<12089> A_IWL<12088> A_IWL<12087> A_IWL<12086> A_IWL<12085> A_IWL<12084> A_IWL<12083> A_IWL<12082> A_IWL<12081> A_IWL<12080> A_IWL<12079> A_IWL<12078> A_IWL<12077> A_IWL<12076> A_IWL<12075> A_IWL<12074> A_IWL<12073> A_IWL<12072> A_IWL<12071> A_IWL<12070> A_IWL<12069> A_IWL<12068> A_IWL<12067> A_IWL<12066> A_IWL<12065> A_IWL<12064> A_IWL<12063> A_IWL<12062> A_IWL<12061> A_IWL<12060> A_IWL<12059> A_IWL<12058> A_IWL<12057> A_IWL<12056> A_IWL<12055> A_IWL<12054> A_IWL<12053> A_IWL<12052> A_IWL<12051> A_IWL<12050> A_IWL<12049> A_IWL<12048> A_IWL<12047> A_IWL<12046> A_IWL<12045> A_IWL<12044> A_IWL<12043> A_IWL<12042> A_IWL<12041> A_IWL<12040> A_IWL<12039> A_IWL<12038> A_IWL<12037> A_IWL<12036> A_IWL<12035> A_IWL<12034> A_IWL<12033> A_IWL<12032> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<46> A_BLC<93> A_BLC<92> A_BLC_TOP<93> A_BLC_TOP<92> A_BLT<93> A_BLT<92> A_BLT_TOP<93> A_BLT_TOP<92> A_IWL<11775> A_IWL<11774> A_IWL<11773> A_IWL<11772> A_IWL<11771> A_IWL<11770> A_IWL<11769> A_IWL<11768> A_IWL<11767> A_IWL<11766> A_IWL<11765> A_IWL<11764> A_IWL<11763> A_IWL<11762> A_IWL<11761> A_IWL<11760> A_IWL<11759> A_IWL<11758> A_IWL<11757> A_IWL<11756> A_IWL<11755> A_IWL<11754> A_IWL<11753> A_IWL<11752> A_IWL<11751> A_IWL<11750> A_IWL<11749> A_IWL<11748> A_IWL<11747> A_IWL<11746> A_IWL<11745> A_IWL<11744> A_IWL<11743> A_IWL<11742> A_IWL<11741> A_IWL<11740> A_IWL<11739> A_IWL<11738> A_IWL<11737> A_IWL<11736> A_IWL<11735> A_IWL<11734> A_IWL<11733> A_IWL<11732> A_IWL<11731> A_IWL<11730> A_IWL<11729> A_IWL<11728> A_IWL<11727> A_IWL<11726> A_IWL<11725> A_IWL<11724> A_IWL<11723> A_IWL<11722> A_IWL<11721> A_IWL<11720> A_IWL<11719> A_IWL<11718> A_IWL<11717> A_IWL<11716> A_IWL<11715> A_IWL<11714> A_IWL<11713> A_IWL<11712> A_IWL<11711> A_IWL<11710> A_IWL<11709> A_IWL<11708> A_IWL<11707> A_IWL<11706> A_IWL<11705> A_IWL<11704> A_IWL<11703> A_IWL<11702> A_IWL<11701> A_IWL<11700> A_IWL<11699> A_IWL<11698> A_IWL<11697> A_IWL<11696> A_IWL<11695> A_IWL<11694> A_IWL<11693> A_IWL<11692> A_IWL<11691> A_IWL<11690> A_IWL<11689> A_IWL<11688> A_IWL<11687> A_IWL<11686> A_IWL<11685> A_IWL<11684> A_IWL<11683> A_IWL<11682> A_IWL<11681> A_IWL<11680> A_IWL<11679> A_IWL<11678> A_IWL<11677> A_IWL<11676> A_IWL<11675> A_IWL<11674> A_IWL<11673> A_IWL<11672> A_IWL<11671> A_IWL<11670> A_IWL<11669> A_IWL<11668> A_IWL<11667> A_IWL<11666> A_IWL<11665> A_IWL<11664> A_IWL<11663> A_IWL<11662> A_IWL<11661> A_IWL<11660> A_IWL<11659> A_IWL<11658> A_IWL<11657> A_IWL<11656> A_IWL<11655> A_IWL<11654> A_IWL<11653> A_IWL<11652> A_IWL<11651> A_IWL<11650> A_IWL<11649> A_IWL<11648> A_IWL<11647> A_IWL<11646> A_IWL<11645> A_IWL<11644> A_IWL<11643> A_IWL<11642> A_IWL<11641> A_IWL<11640> A_IWL<11639> A_IWL<11638> A_IWL<11637> A_IWL<11636> A_IWL<11635> A_IWL<11634> A_IWL<11633> A_IWL<11632> A_IWL<11631> A_IWL<11630> A_IWL<11629> A_IWL<11628> A_IWL<11627> A_IWL<11626> A_IWL<11625> A_IWL<11624> A_IWL<11623> A_IWL<11622> A_IWL<11621> A_IWL<11620> A_IWL<11619> A_IWL<11618> A_IWL<11617> A_IWL<11616> A_IWL<11615> A_IWL<11614> A_IWL<11613> A_IWL<11612> A_IWL<11611> A_IWL<11610> A_IWL<11609> A_IWL<11608> A_IWL<11607> A_IWL<11606> A_IWL<11605> A_IWL<11604> A_IWL<11603> A_IWL<11602> A_IWL<11601> A_IWL<11600> A_IWL<11599> A_IWL<11598> A_IWL<11597> A_IWL<11596> A_IWL<11595> A_IWL<11594> A_IWL<11593> A_IWL<11592> A_IWL<11591> A_IWL<11590> A_IWL<11589> A_IWL<11588> A_IWL<11587> A_IWL<11586> A_IWL<11585> A_IWL<11584> A_IWL<11583> A_IWL<11582> A_IWL<11581> A_IWL<11580> A_IWL<11579> A_IWL<11578> A_IWL<11577> A_IWL<11576> A_IWL<11575> A_IWL<11574> A_IWL<11573> A_IWL<11572> A_IWL<11571> A_IWL<11570> A_IWL<11569> A_IWL<11568> A_IWL<11567> A_IWL<11566> A_IWL<11565> A_IWL<11564> A_IWL<11563> A_IWL<11562> A_IWL<11561> A_IWL<11560> A_IWL<11559> A_IWL<11558> A_IWL<11557> A_IWL<11556> A_IWL<11555> A_IWL<11554> A_IWL<11553> A_IWL<11552> A_IWL<11551> A_IWL<11550> A_IWL<11549> A_IWL<11548> A_IWL<11547> A_IWL<11546> A_IWL<11545> A_IWL<11544> A_IWL<11543> A_IWL<11542> A_IWL<11541> A_IWL<11540> A_IWL<11539> A_IWL<11538> A_IWL<11537> A_IWL<11536> A_IWL<11535> A_IWL<11534> A_IWL<11533> A_IWL<11532> A_IWL<11531> A_IWL<11530> A_IWL<11529> A_IWL<11528> A_IWL<11527> A_IWL<11526> A_IWL<11525> A_IWL<11524> A_IWL<11523> A_IWL<11522> A_IWL<11521> A_IWL<11520> A_IWL<12031> A_IWL<12030> A_IWL<12029> A_IWL<12028> A_IWL<12027> A_IWL<12026> A_IWL<12025> A_IWL<12024> A_IWL<12023> A_IWL<12022> A_IWL<12021> A_IWL<12020> A_IWL<12019> A_IWL<12018> A_IWL<12017> A_IWL<12016> A_IWL<12015> A_IWL<12014> A_IWL<12013> A_IWL<12012> A_IWL<12011> A_IWL<12010> A_IWL<12009> A_IWL<12008> A_IWL<12007> A_IWL<12006> A_IWL<12005> A_IWL<12004> A_IWL<12003> A_IWL<12002> A_IWL<12001> A_IWL<12000> A_IWL<11999> A_IWL<11998> A_IWL<11997> A_IWL<11996> A_IWL<11995> A_IWL<11994> A_IWL<11993> A_IWL<11992> A_IWL<11991> A_IWL<11990> A_IWL<11989> A_IWL<11988> A_IWL<11987> A_IWL<11986> A_IWL<11985> A_IWL<11984> A_IWL<11983> A_IWL<11982> A_IWL<11981> A_IWL<11980> A_IWL<11979> A_IWL<11978> A_IWL<11977> A_IWL<11976> A_IWL<11975> A_IWL<11974> A_IWL<11973> A_IWL<11972> A_IWL<11971> A_IWL<11970> A_IWL<11969> A_IWL<11968> A_IWL<11967> A_IWL<11966> A_IWL<11965> A_IWL<11964> A_IWL<11963> A_IWL<11962> A_IWL<11961> A_IWL<11960> A_IWL<11959> A_IWL<11958> A_IWL<11957> A_IWL<11956> A_IWL<11955> A_IWL<11954> A_IWL<11953> A_IWL<11952> A_IWL<11951> A_IWL<11950> A_IWL<11949> A_IWL<11948> A_IWL<11947> A_IWL<11946> A_IWL<11945> A_IWL<11944> A_IWL<11943> A_IWL<11942> A_IWL<11941> A_IWL<11940> A_IWL<11939> A_IWL<11938> A_IWL<11937> A_IWL<11936> A_IWL<11935> A_IWL<11934> A_IWL<11933> A_IWL<11932> A_IWL<11931> A_IWL<11930> A_IWL<11929> A_IWL<11928> A_IWL<11927> A_IWL<11926> A_IWL<11925> A_IWL<11924> A_IWL<11923> A_IWL<11922> A_IWL<11921> A_IWL<11920> A_IWL<11919> A_IWL<11918> A_IWL<11917> A_IWL<11916> A_IWL<11915> A_IWL<11914> A_IWL<11913> A_IWL<11912> A_IWL<11911> A_IWL<11910> A_IWL<11909> A_IWL<11908> A_IWL<11907> A_IWL<11906> A_IWL<11905> A_IWL<11904> A_IWL<11903> A_IWL<11902> A_IWL<11901> A_IWL<11900> A_IWL<11899> A_IWL<11898> A_IWL<11897> A_IWL<11896> A_IWL<11895> A_IWL<11894> A_IWL<11893> A_IWL<11892> A_IWL<11891> A_IWL<11890> A_IWL<11889> A_IWL<11888> A_IWL<11887> A_IWL<11886> A_IWL<11885> A_IWL<11884> A_IWL<11883> A_IWL<11882> A_IWL<11881> A_IWL<11880> A_IWL<11879> A_IWL<11878> A_IWL<11877> A_IWL<11876> A_IWL<11875> A_IWL<11874> A_IWL<11873> A_IWL<11872> A_IWL<11871> A_IWL<11870> A_IWL<11869> A_IWL<11868> A_IWL<11867> A_IWL<11866> A_IWL<11865> A_IWL<11864> A_IWL<11863> A_IWL<11862> A_IWL<11861> A_IWL<11860> A_IWL<11859> A_IWL<11858> A_IWL<11857> A_IWL<11856> A_IWL<11855> A_IWL<11854> A_IWL<11853> A_IWL<11852> A_IWL<11851> A_IWL<11850> A_IWL<11849> A_IWL<11848> A_IWL<11847> A_IWL<11846> A_IWL<11845> A_IWL<11844> A_IWL<11843> A_IWL<11842> A_IWL<11841> A_IWL<11840> A_IWL<11839> A_IWL<11838> A_IWL<11837> A_IWL<11836> A_IWL<11835> A_IWL<11834> A_IWL<11833> A_IWL<11832> A_IWL<11831> A_IWL<11830> A_IWL<11829> A_IWL<11828> A_IWL<11827> A_IWL<11826> A_IWL<11825> A_IWL<11824> A_IWL<11823> A_IWL<11822> A_IWL<11821> A_IWL<11820> A_IWL<11819> A_IWL<11818> A_IWL<11817> A_IWL<11816> A_IWL<11815> A_IWL<11814> A_IWL<11813> A_IWL<11812> A_IWL<11811> A_IWL<11810> A_IWL<11809> A_IWL<11808> A_IWL<11807> A_IWL<11806> A_IWL<11805> A_IWL<11804> A_IWL<11803> A_IWL<11802> A_IWL<11801> A_IWL<11800> A_IWL<11799> A_IWL<11798> A_IWL<11797> A_IWL<11796> A_IWL<11795> A_IWL<11794> A_IWL<11793> A_IWL<11792> A_IWL<11791> A_IWL<11790> A_IWL<11789> A_IWL<11788> A_IWL<11787> A_IWL<11786> A_IWL<11785> A_IWL<11784> A_IWL<11783> A_IWL<11782> A_IWL<11781> A_IWL<11780> A_IWL<11779> A_IWL<11778> A_IWL<11777> A_IWL<11776> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<45> A_BLC<91> A_BLC<90> A_BLC_TOP<91> A_BLC_TOP<90> A_BLT<91> A_BLT<90> A_BLT_TOP<91> A_BLT_TOP<90> A_IWL<11519> A_IWL<11518> A_IWL<11517> A_IWL<11516> A_IWL<11515> A_IWL<11514> A_IWL<11513> A_IWL<11512> A_IWL<11511> A_IWL<11510> A_IWL<11509> A_IWL<11508> A_IWL<11507> A_IWL<11506> A_IWL<11505> A_IWL<11504> A_IWL<11503> A_IWL<11502> A_IWL<11501> A_IWL<11500> A_IWL<11499> A_IWL<11498> A_IWL<11497> A_IWL<11496> A_IWL<11495> A_IWL<11494> A_IWL<11493> A_IWL<11492> A_IWL<11491> A_IWL<11490> A_IWL<11489> A_IWL<11488> A_IWL<11487> A_IWL<11486> A_IWL<11485> A_IWL<11484> A_IWL<11483> A_IWL<11482> A_IWL<11481> A_IWL<11480> A_IWL<11479> A_IWL<11478> A_IWL<11477> A_IWL<11476> A_IWL<11475> A_IWL<11474> A_IWL<11473> A_IWL<11472> A_IWL<11471> A_IWL<11470> A_IWL<11469> A_IWL<11468> A_IWL<11467> A_IWL<11466> A_IWL<11465> A_IWL<11464> A_IWL<11463> A_IWL<11462> A_IWL<11461> A_IWL<11460> A_IWL<11459> A_IWL<11458> A_IWL<11457> A_IWL<11456> A_IWL<11455> A_IWL<11454> A_IWL<11453> A_IWL<11452> A_IWL<11451> A_IWL<11450> A_IWL<11449> A_IWL<11448> A_IWL<11447> A_IWL<11446> A_IWL<11445> A_IWL<11444> A_IWL<11443> A_IWL<11442> A_IWL<11441> A_IWL<11440> A_IWL<11439> A_IWL<11438> A_IWL<11437> A_IWL<11436> A_IWL<11435> A_IWL<11434> A_IWL<11433> A_IWL<11432> A_IWL<11431> A_IWL<11430> A_IWL<11429> A_IWL<11428> A_IWL<11427> A_IWL<11426> A_IWL<11425> A_IWL<11424> A_IWL<11423> A_IWL<11422> A_IWL<11421> A_IWL<11420> A_IWL<11419> A_IWL<11418> A_IWL<11417> A_IWL<11416> A_IWL<11415> A_IWL<11414> A_IWL<11413> A_IWL<11412> A_IWL<11411> A_IWL<11410> A_IWL<11409> A_IWL<11408> A_IWL<11407> A_IWL<11406> A_IWL<11405> A_IWL<11404> A_IWL<11403> A_IWL<11402> A_IWL<11401> A_IWL<11400> A_IWL<11399> A_IWL<11398> A_IWL<11397> A_IWL<11396> A_IWL<11395> A_IWL<11394> A_IWL<11393> A_IWL<11392> A_IWL<11391> A_IWL<11390> A_IWL<11389> A_IWL<11388> A_IWL<11387> A_IWL<11386> A_IWL<11385> A_IWL<11384> A_IWL<11383> A_IWL<11382> A_IWL<11381> A_IWL<11380> A_IWL<11379> A_IWL<11378> A_IWL<11377> A_IWL<11376> A_IWL<11375> A_IWL<11374> A_IWL<11373> A_IWL<11372> A_IWL<11371> A_IWL<11370> A_IWL<11369> A_IWL<11368> A_IWL<11367> A_IWL<11366> A_IWL<11365> A_IWL<11364> A_IWL<11363> A_IWL<11362> A_IWL<11361> A_IWL<11360> A_IWL<11359> A_IWL<11358> A_IWL<11357> A_IWL<11356> A_IWL<11355> A_IWL<11354> A_IWL<11353> A_IWL<11352> A_IWL<11351> A_IWL<11350> A_IWL<11349> A_IWL<11348> A_IWL<11347> A_IWL<11346> A_IWL<11345> A_IWL<11344> A_IWL<11343> A_IWL<11342> A_IWL<11341> A_IWL<11340> A_IWL<11339> A_IWL<11338> A_IWL<11337> A_IWL<11336> A_IWL<11335> A_IWL<11334> A_IWL<11333> A_IWL<11332> A_IWL<11331> A_IWL<11330> A_IWL<11329> A_IWL<11328> A_IWL<11327> A_IWL<11326> A_IWL<11325> A_IWL<11324> A_IWL<11323> A_IWL<11322> A_IWL<11321> A_IWL<11320> A_IWL<11319> A_IWL<11318> A_IWL<11317> A_IWL<11316> A_IWL<11315> A_IWL<11314> A_IWL<11313> A_IWL<11312> A_IWL<11311> A_IWL<11310> A_IWL<11309> A_IWL<11308> A_IWL<11307> A_IWL<11306> A_IWL<11305> A_IWL<11304> A_IWL<11303> A_IWL<11302> A_IWL<11301> A_IWL<11300> A_IWL<11299> A_IWL<11298> A_IWL<11297> A_IWL<11296> A_IWL<11295> A_IWL<11294> A_IWL<11293> A_IWL<11292> A_IWL<11291> A_IWL<11290> A_IWL<11289> A_IWL<11288> A_IWL<11287> A_IWL<11286> A_IWL<11285> A_IWL<11284> A_IWL<11283> A_IWL<11282> A_IWL<11281> A_IWL<11280> A_IWL<11279> A_IWL<11278> A_IWL<11277> A_IWL<11276> A_IWL<11275> A_IWL<11274> A_IWL<11273> A_IWL<11272> A_IWL<11271> A_IWL<11270> A_IWL<11269> A_IWL<11268> A_IWL<11267> A_IWL<11266> A_IWL<11265> A_IWL<11264> A_IWL<11775> A_IWL<11774> A_IWL<11773> A_IWL<11772> A_IWL<11771> A_IWL<11770> A_IWL<11769> A_IWL<11768> A_IWL<11767> A_IWL<11766> A_IWL<11765> A_IWL<11764> A_IWL<11763> A_IWL<11762> A_IWL<11761> A_IWL<11760> A_IWL<11759> A_IWL<11758> A_IWL<11757> A_IWL<11756> A_IWL<11755> A_IWL<11754> A_IWL<11753> A_IWL<11752> A_IWL<11751> A_IWL<11750> A_IWL<11749> A_IWL<11748> A_IWL<11747> A_IWL<11746> A_IWL<11745> A_IWL<11744> A_IWL<11743> A_IWL<11742> A_IWL<11741> A_IWL<11740> A_IWL<11739> A_IWL<11738> A_IWL<11737> A_IWL<11736> A_IWL<11735> A_IWL<11734> A_IWL<11733> A_IWL<11732> A_IWL<11731> A_IWL<11730> A_IWL<11729> A_IWL<11728> A_IWL<11727> A_IWL<11726> A_IWL<11725> A_IWL<11724> A_IWL<11723> A_IWL<11722> A_IWL<11721> A_IWL<11720> A_IWL<11719> A_IWL<11718> A_IWL<11717> A_IWL<11716> A_IWL<11715> A_IWL<11714> A_IWL<11713> A_IWL<11712> A_IWL<11711> A_IWL<11710> A_IWL<11709> A_IWL<11708> A_IWL<11707> A_IWL<11706> A_IWL<11705> A_IWL<11704> A_IWL<11703> A_IWL<11702> A_IWL<11701> A_IWL<11700> A_IWL<11699> A_IWL<11698> A_IWL<11697> A_IWL<11696> A_IWL<11695> A_IWL<11694> A_IWL<11693> A_IWL<11692> A_IWL<11691> A_IWL<11690> A_IWL<11689> A_IWL<11688> A_IWL<11687> A_IWL<11686> A_IWL<11685> A_IWL<11684> A_IWL<11683> A_IWL<11682> A_IWL<11681> A_IWL<11680> A_IWL<11679> A_IWL<11678> A_IWL<11677> A_IWL<11676> A_IWL<11675> A_IWL<11674> A_IWL<11673> A_IWL<11672> A_IWL<11671> A_IWL<11670> A_IWL<11669> A_IWL<11668> A_IWL<11667> A_IWL<11666> A_IWL<11665> A_IWL<11664> A_IWL<11663> A_IWL<11662> A_IWL<11661> A_IWL<11660> A_IWL<11659> A_IWL<11658> A_IWL<11657> A_IWL<11656> A_IWL<11655> A_IWL<11654> A_IWL<11653> A_IWL<11652> A_IWL<11651> A_IWL<11650> A_IWL<11649> A_IWL<11648> A_IWL<11647> A_IWL<11646> A_IWL<11645> A_IWL<11644> A_IWL<11643> A_IWL<11642> A_IWL<11641> A_IWL<11640> A_IWL<11639> A_IWL<11638> A_IWL<11637> A_IWL<11636> A_IWL<11635> A_IWL<11634> A_IWL<11633> A_IWL<11632> A_IWL<11631> A_IWL<11630> A_IWL<11629> A_IWL<11628> A_IWL<11627> A_IWL<11626> A_IWL<11625> A_IWL<11624> A_IWL<11623> A_IWL<11622> A_IWL<11621> A_IWL<11620> A_IWL<11619> A_IWL<11618> A_IWL<11617> A_IWL<11616> A_IWL<11615> A_IWL<11614> A_IWL<11613> A_IWL<11612> A_IWL<11611> A_IWL<11610> A_IWL<11609> A_IWL<11608> A_IWL<11607> A_IWL<11606> A_IWL<11605> A_IWL<11604> A_IWL<11603> A_IWL<11602> A_IWL<11601> A_IWL<11600> A_IWL<11599> A_IWL<11598> A_IWL<11597> A_IWL<11596> A_IWL<11595> A_IWL<11594> A_IWL<11593> A_IWL<11592> A_IWL<11591> A_IWL<11590> A_IWL<11589> A_IWL<11588> A_IWL<11587> A_IWL<11586> A_IWL<11585> A_IWL<11584> A_IWL<11583> A_IWL<11582> A_IWL<11581> A_IWL<11580> A_IWL<11579> A_IWL<11578> A_IWL<11577> A_IWL<11576> A_IWL<11575> A_IWL<11574> A_IWL<11573> A_IWL<11572> A_IWL<11571> A_IWL<11570> A_IWL<11569> A_IWL<11568> A_IWL<11567> A_IWL<11566> A_IWL<11565> A_IWL<11564> A_IWL<11563> A_IWL<11562> A_IWL<11561> A_IWL<11560> A_IWL<11559> A_IWL<11558> A_IWL<11557> A_IWL<11556> A_IWL<11555> A_IWL<11554> A_IWL<11553> A_IWL<11552> A_IWL<11551> A_IWL<11550> A_IWL<11549> A_IWL<11548> A_IWL<11547> A_IWL<11546> A_IWL<11545> A_IWL<11544> A_IWL<11543> A_IWL<11542> A_IWL<11541> A_IWL<11540> A_IWL<11539> A_IWL<11538> A_IWL<11537> A_IWL<11536> A_IWL<11535> A_IWL<11534> A_IWL<11533> A_IWL<11532> A_IWL<11531> A_IWL<11530> A_IWL<11529> A_IWL<11528> A_IWL<11527> A_IWL<11526> A_IWL<11525> A_IWL<11524> A_IWL<11523> A_IWL<11522> A_IWL<11521> A_IWL<11520> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<44> A_BLC<89> A_BLC<88> A_BLC_TOP<89> A_BLC_TOP<88> A_BLT<89> A_BLT<88> A_BLT_TOP<89> A_BLT_TOP<88> A_IWL<11263> A_IWL<11262> A_IWL<11261> A_IWL<11260> A_IWL<11259> A_IWL<11258> A_IWL<11257> A_IWL<11256> A_IWL<11255> A_IWL<11254> A_IWL<11253> A_IWL<11252> A_IWL<11251> A_IWL<11250> A_IWL<11249> A_IWL<11248> A_IWL<11247> A_IWL<11246> A_IWL<11245> A_IWL<11244> A_IWL<11243> A_IWL<11242> A_IWL<11241> A_IWL<11240> A_IWL<11239> A_IWL<11238> A_IWL<11237> A_IWL<11236> A_IWL<11235> A_IWL<11234> A_IWL<11233> A_IWL<11232> A_IWL<11231> A_IWL<11230> A_IWL<11229> A_IWL<11228> A_IWL<11227> A_IWL<11226> A_IWL<11225> A_IWL<11224> A_IWL<11223> A_IWL<11222> A_IWL<11221> A_IWL<11220> A_IWL<11219> A_IWL<11218> A_IWL<11217> A_IWL<11216> A_IWL<11215> A_IWL<11214> A_IWL<11213> A_IWL<11212> A_IWL<11211> A_IWL<11210> A_IWL<11209> A_IWL<11208> A_IWL<11207> A_IWL<11206> A_IWL<11205> A_IWL<11204> A_IWL<11203> A_IWL<11202> A_IWL<11201> A_IWL<11200> A_IWL<11199> A_IWL<11198> A_IWL<11197> A_IWL<11196> A_IWL<11195> A_IWL<11194> A_IWL<11193> A_IWL<11192> A_IWL<11191> A_IWL<11190> A_IWL<11189> A_IWL<11188> A_IWL<11187> A_IWL<11186> A_IWL<11185> A_IWL<11184> A_IWL<11183> A_IWL<11182> A_IWL<11181> A_IWL<11180> A_IWL<11179> A_IWL<11178> A_IWL<11177> A_IWL<11176> A_IWL<11175> A_IWL<11174> A_IWL<11173> A_IWL<11172> A_IWL<11171> A_IWL<11170> A_IWL<11169> A_IWL<11168> A_IWL<11167> A_IWL<11166> A_IWL<11165> A_IWL<11164> A_IWL<11163> A_IWL<11162> A_IWL<11161> A_IWL<11160> A_IWL<11159> A_IWL<11158> A_IWL<11157> A_IWL<11156> A_IWL<11155> A_IWL<11154> A_IWL<11153> A_IWL<11152> A_IWL<11151> A_IWL<11150> A_IWL<11149> A_IWL<11148> A_IWL<11147> A_IWL<11146> A_IWL<11145> A_IWL<11144> A_IWL<11143> A_IWL<11142> A_IWL<11141> A_IWL<11140> A_IWL<11139> A_IWL<11138> A_IWL<11137> A_IWL<11136> A_IWL<11135> A_IWL<11134> A_IWL<11133> A_IWL<11132> A_IWL<11131> A_IWL<11130> A_IWL<11129> A_IWL<11128> A_IWL<11127> A_IWL<11126> A_IWL<11125> A_IWL<11124> A_IWL<11123> A_IWL<11122> A_IWL<11121> A_IWL<11120> A_IWL<11119> A_IWL<11118> A_IWL<11117> A_IWL<11116> A_IWL<11115> A_IWL<11114> A_IWL<11113> A_IWL<11112> A_IWL<11111> A_IWL<11110> A_IWL<11109> A_IWL<11108> A_IWL<11107> A_IWL<11106> A_IWL<11105> A_IWL<11104> A_IWL<11103> A_IWL<11102> A_IWL<11101> A_IWL<11100> A_IWL<11099> A_IWL<11098> A_IWL<11097> A_IWL<11096> A_IWL<11095> A_IWL<11094> A_IWL<11093> A_IWL<11092> A_IWL<11091> A_IWL<11090> A_IWL<11089> A_IWL<11088> A_IWL<11087> A_IWL<11086> A_IWL<11085> A_IWL<11084> A_IWL<11083> A_IWL<11082> A_IWL<11081> A_IWL<11080> A_IWL<11079> A_IWL<11078> A_IWL<11077> A_IWL<11076> A_IWL<11075> A_IWL<11074> A_IWL<11073> A_IWL<11072> A_IWL<11071> A_IWL<11070> A_IWL<11069> A_IWL<11068> A_IWL<11067> A_IWL<11066> A_IWL<11065> A_IWL<11064> A_IWL<11063> A_IWL<11062> A_IWL<11061> A_IWL<11060> A_IWL<11059> A_IWL<11058> A_IWL<11057> A_IWL<11056> A_IWL<11055> A_IWL<11054> A_IWL<11053> A_IWL<11052> A_IWL<11051> A_IWL<11050> A_IWL<11049> A_IWL<11048> A_IWL<11047> A_IWL<11046> A_IWL<11045> A_IWL<11044> A_IWL<11043> A_IWL<11042> A_IWL<11041> A_IWL<11040> A_IWL<11039> A_IWL<11038> A_IWL<11037> A_IWL<11036> A_IWL<11035> A_IWL<11034> A_IWL<11033> A_IWL<11032> A_IWL<11031> A_IWL<11030> A_IWL<11029> A_IWL<11028> A_IWL<11027> A_IWL<11026> A_IWL<11025> A_IWL<11024> A_IWL<11023> A_IWL<11022> A_IWL<11021> A_IWL<11020> A_IWL<11019> A_IWL<11018> A_IWL<11017> A_IWL<11016> A_IWL<11015> A_IWL<11014> A_IWL<11013> A_IWL<11012> A_IWL<11011> A_IWL<11010> A_IWL<11009> A_IWL<11008> A_IWL<11519> A_IWL<11518> A_IWL<11517> A_IWL<11516> A_IWL<11515> A_IWL<11514> A_IWL<11513> A_IWL<11512> A_IWL<11511> A_IWL<11510> A_IWL<11509> A_IWL<11508> A_IWL<11507> A_IWL<11506> A_IWL<11505> A_IWL<11504> A_IWL<11503> A_IWL<11502> A_IWL<11501> A_IWL<11500> A_IWL<11499> A_IWL<11498> A_IWL<11497> A_IWL<11496> A_IWL<11495> A_IWL<11494> A_IWL<11493> A_IWL<11492> A_IWL<11491> A_IWL<11490> A_IWL<11489> A_IWL<11488> A_IWL<11487> A_IWL<11486> A_IWL<11485> A_IWL<11484> A_IWL<11483> A_IWL<11482> A_IWL<11481> A_IWL<11480> A_IWL<11479> A_IWL<11478> A_IWL<11477> A_IWL<11476> A_IWL<11475> A_IWL<11474> A_IWL<11473> A_IWL<11472> A_IWL<11471> A_IWL<11470> A_IWL<11469> A_IWL<11468> A_IWL<11467> A_IWL<11466> A_IWL<11465> A_IWL<11464> A_IWL<11463> A_IWL<11462> A_IWL<11461> A_IWL<11460> A_IWL<11459> A_IWL<11458> A_IWL<11457> A_IWL<11456> A_IWL<11455> A_IWL<11454> A_IWL<11453> A_IWL<11452> A_IWL<11451> A_IWL<11450> A_IWL<11449> A_IWL<11448> A_IWL<11447> A_IWL<11446> A_IWL<11445> A_IWL<11444> A_IWL<11443> A_IWL<11442> A_IWL<11441> A_IWL<11440> A_IWL<11439> A_IWL<11438> A_IWL<11437> A_IWL<11436> A_IWL<11435> A_IWL<11434> A_IWL<11433> A_IWL<11432> A_IWL<11431> A_IWL<11430> A_IWL<11429> A_IWL<11428> A_IWL<11427> A_IWL<11426> A_IWL<11425> A_IWL<11424> A_IWL<11423> A_IWL<11422> A_IWL<11421> A_IWL<11420> A_IWL<11419> A_IWL<11418> A_IWL<11417> A_IWL<11416> A_IWL<11415> A_IWL<11414> A_IWL<11413> A_IWL<11412> A_IWL<11411> A_IWL<11410> A_IWL<11409> A_IWL<11408> A_IWL<11407> A_IWL<11406> A_IWL<11405> A_IWL<11404> A_IWL<11403> A_IWL<11402> A_IWL<11401> A_IWL<11400> A_IWL<11399> A_IWL<11398> A_IWL<11397> A_IWL<11396> A_IWL<11395> A_IWL<11394> A_IWL<11393> A_IWL<11392> A_IWL<11391> A_IWL<11390> A_IWL<11389> A_IWL<11388> A_IWL<11387> A_IWL<11386> A_IWL<11385> A_IWL<11384> A_IWL<11383> A_IWL<11382> A_IWL<11381> A_IWL<11380> A_IWL<11379> A_IWL<11378> A_IWL<11377> A_IWL<11376> A_IWL<11375> A_IWL<11374> A_IWL<11373> A_IWL<11372> A_IWL<11371> A_IWL<11370> A_IWL<11369> A_IWL<11368> A_IWL<11367> A_IWL<11366> A_IWL<11365> A_IWL<11364> A_IWL<11363> A_IWL<11362> A_IWL<11361> A_IWL<11360> A_IWL<11359> A_IWL<11358> A_IWL<11357> A_IWL<11356> A_IWL<11355> A_IWL<11354> A_IWL<11353> A_IWL<11352> A_IWL<11351> A_IWL<11350> A_IWL<11349> A_IWL<11348> A_IWL<11347> A_IWL<11346> A_IWL<11345> A_IWL<11344> A_IWL<11343> A_IWL<11342> A_IWL<11341> A_IWL<11340> A_IWL<11339> A_IWL<11338> A_IWL<11337> A_IWL<11336> A_IWL<11335> A_IWL<11334> A_IWL<11333> A_IWL<11332> A_IWL<11331> A_IWL<11330> A_IWL<11329> A_IWL<11328> A_IWL<11327> A_IWL<11326> A_IWL<11325> A_IWL<11324> A_IWL<11323> A_IWL<11322> A_IWL<11321> A_IWL<11320> A_IWL<11319> A_IWL<11318> A_IWL<11317> A_IWL<11316> A_IWL<11315> A_IWL<11314> A_IWL<11313> A_IWL<11312> A_IWL<11311> A_IWL<11310> A_IWL<11309> A_IWL<11308> A_IWL<11307> A_IWL<11306> A_IWL<11305> A_IWL<11304> A_IWL<11303> A_IWL<11302> A_IWL<11301> A_IWL<11300> A_IWL<11299> A_IWL<11298> A_IWL<11297> A_IWL<11296> A_IWL<11295> A_IWL<11294> A_IWL<11293> A_IWL<11292> A_IWL<11291> A_IWL<11290> A_IWL<11289> A_IWL<11288> A_IWL<11287> A_IWL<11286> A_IWL<11285> A_IWL<11284> A_IWL<11283> A_IWL<11282> A_IWL<11281> A_IWL<11280> A_IWL<11279> A_IWL<11278> A_IWL<11277> A_IWL<11276> A_IWL<11275> A_IWL<11274> A_IWL<11273> A_IWL<11272> A_IWL<11271> A_IWL<11270> A_IWL<11269> A_IWL<11268> A_IWL<11267> A_IWL<11266> A_IWL<11265> A_IWL<11264> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<43> A_BLC<87> A_BLC<86> A_BLC_TOP<87> A_BLC_TOP<86> A_BLT<87> A_BLT<86> A_BLT_TOP<87> A_BLT_TOP<86> A_IWL<11007> A_IWL<11006> A_IWL<11005> A_IWL<11004> A_IWL<11003> A_IWL<11002> A_IWL<11001> A_IWL<11000> A_IWL<10999> A_IWL<10998> A_IWL<10997> A_IWL<10996> A_IWL<10995> A_IWL<10994> A_IWL<10993> A_IWL<10992> A_IWL<10991> A_IWL<10990> A_IWL<10989> A_IWL<10988> A_IWL<10987> A_IWL<10986> A_IWL<10985> A_IWL<10984> A_IWL<10983> A_IWL<10982> A_IWL<10981> A_IWL<10980> A_IWL<10979> A_IWL<10978> A_IWL<10977> A_IWL<10976> A_IWL<10975> A_IWL<10974> A_IWL<10973> A_IWL<10972> A_IWL<10971> A_IWL<10970> A_IWL<10969> A_IWL<10968> A_IWL<10967> A_IWL<10966> A_IWL<10965> A_IWL<10964> A_IWL<10963> A_IWL<10962> A_IWL<10961> A_IWL<10960> A_IWL<10959> A_IWL<10958> A_IWL<10957> A_IWL<10956> A_IWL<10955> A_IWL<10954> A_IWL<10953> A_IWL<10952> A_IWL<10951> A_IWL<10950> A_IWL<10949> A_IWL<10948> A_IWL<10947> A_IWL<10946> A_IWL<10945> A_IWL<10944> A_IWL<10943> A_IWL<10942> A_IWL<10941> A_IWL<10940> A_IWL<10939> A_IWL<10938> A_IWL<10937> A_IWL<10936> A_IWL<10935> A_IWL<10934> A_IWL<10933> A_IWL<10932> A_IWL<10931> A_IWL<10930> A_IWL<10929> A_IWL<10928> A_IWL<10927> A_IWL<10926> A_IWL<10925> A_IWL<10924> A_IWL<10923> A_IWL<10922> A_IWL<10921> A_IWL<10920> A_IWL<10919> A_IWL<10918> A_IWL<10917> A_IWL<10916> A_IWL<10915> A_IWL<10914> A_IWL<10913> A_IWL<10912> A_IWL<10911> A_IWL<10910> A_IWL<10909> A_IWL<10908> A_IWL<10907> A_IWL<10906> A_IWL<10905> A_IWL<10904> A_IWL<10903> A_IWL<10902> A_IWL<10901> A_IWL<10900> A_IWL<10899> A_IWL<10898> A_IWL<10897> A_IWL<10896> A_IWL<10895> A_IWL<10894> A_IWL<10893> A_IWL<10892> A_IWL<10891> A_IWL<10890> A_IWL<10889> A_IWL<10888> A_IWL<10887> A_IWL<10886> A_IWL<10885> A_IWL<10884> A_IWL<10883> A_IWL<10882> A_IWL<10881> A_IWL<10880> A_IWL<10879> A_IWL<10878> A_IWL<10877> A_IWL<10876> A_IWL<10875> A_IWL<10874> A_IWL<10873> A_IWL<10872> A_IWL<10871> A_IWL<10870> A_IWL<10869> A_IWL<10868> A_IWL<10867> A_IWL<10866> A_IWL<10865> A_IWL<10864> A_IWL<10863> A_IWL<10862> A_IWL<10861> A_IWL<10860> A_IWL<10859> A_IWL<10858> A_IWL<10857> A_IWL<10856> A_IWL<10855> A_IWL<10854> A_IWL<10853> A_IWL<10852> A_IWL<10851> A_IWL<10850> A_IWL<10849> A_IWL<10848> A_IWL<10847> A_IWL<10846> A_IWL<10845> A_IWL<10844> A_IWL<10843> A_IWL<10842> A_IWL<10841> A_IWL<10840> A_IWL<10839> A_IWL<10838> A_IWL<10837> A_IWL<10836> A_IWL<10835> A_IWL<10834> A_IWL<10833> A_IWL<10832> A_IWL<10831> A_IWL<10830> A_IWL<10829> A_IWL<10828> A_IWL<10827> A_IWL<10826> A_IWL<10825> A_IWL<10824> A_IWL<10823> A_IWL<10822> A_IWL<10821> A_IWL<10820> A_IWL<10819> A_IWL<10818> A_IWL<10817> A_IWL<10816> A_IWL<10815> A_IWL<10814> A_IWL<10813> A_IWL<10812> A_IWL<10811> A_IWL<10810> A_IWL<10809> A_IWL<10808> A_IWL<10807> A_IWL<10806> A_IWL<10805> A_IWL<10804> A_IWL<10803> A_IWL<10802> A_IWL<10801> A_IWL<10800> A_IWL<10799> A_IWL<10798> A_IWL<10797> A_IWL<10796> A_IWL<10795> A_IWL<10794> A_IWL<10793> A_IWL<10792> A_IWL<10791> A_IWL<10790> A_IWL<10789> A_IWL<10788> A_IWL<10787> A_IWL<10786> A_IWL<10785> A_IWL<10784> A_IWL<10783> A_IWL<10782> A_IWL<10781> A_IWL<10780> A_IWL<10779> A_IWL<10778> A_IWL<10777> A_IWL<10776> A_IWL<10775> A_IWL<10774> A_IWL<10773> A_IWL<10772> A_IWL<10771> A_IWL<10770> A_IWL<10769> A_IWL<10768> A_IWL<10767> A_IWL<10766> A_IWL<10765> A_IWL<10764> A_IWL<10763> A_IWL<10762> A_IWL<10761> A_IWL<10760> A_IWL<10759> A_IWL<10758> A_IWL<10757> A_IWL<10756> A_IWL<10755> A_IWL<10754> A_IWL<10753> A_IWL<10752> A_IWL<11263> A_IWL<11262> A_IWL<11261> A_IWL<11260> A_IWL<11259> A_IWL<11258> A_IWL<11257> A_IWL<11256> A_IWL<11255> A_IWL<11254> A_IWL<11253> A_IWL<11252> A_IWL<11251> A_IWL<11250> A_IWL<11249> A_IWL<11248> A_IWL<11247> A_IWL<11246> A_IWL<11245> A_IWL<11244> A_IWL<11243> A_IWL<11242> A_IWL<11241> A_IWL<11240> A_IWL<11239> A_IWL<11238> A_IWL<11237> A_IWL<11236> A_IWL<11235> A_IWL<11234> A_IWL<11233> A_IWL<11232> A_IWL<11231> A_IWL<11230> A_IWL<11229> A_IWL<11228> A_IWL<11227> A_IWL<11226> A_IWL<11225> A_IWL<11224> A_IWL<11223> A_IWL<11222> A_IWL<11221> A_IWL<11220> A_IWL<11219> A_IWL<11218> A_IWL<11217> A_IWL<11216> A_IWL<11215> A_IWL<11214> A_IWL<11213> A_IWL<11212> A_IWL<11211> A_IWL<11210> A_IWL<11209> A_IWL<11208> A_IWL<11207> A_IWL<11206> A_IWL<11205> A_IWL<11204> A_IWL<11203> A_IWL<11202> A_IWL<11201> A_IWL<11200> A_IWL<11199> A_IWL<11198> A_IWL<11197> A_IWL<11196> A_IWL<11195> A_IWL<11194> A_IWL<11193> A_IWL<11192> A_IWL<11191> A_IWL<11190> A_IWL<11189> A_IWL<11188> A_IWL<11187> A_IWL<11186> A_IWL<11185> A_IWL<11184> A_IWL<11183> A_IWL<11182> A_IWL<11181> A_IWL<11180> A_IWL<11179> A_IWL<11178> A_IWL<11177> A_IWL<11176> A_IWL<11175> A_IWL<11174> A_IWL<11173> A_IWL<11172> A_IWL<11171> A_IWL<11170> A_IWL<11169> A_IWL<11168> A_IWL<11167> A_IWL<11166> A_IWL<11165> A_IWL<11164> A_IWL<11163> A_IWL<11162> A_IWL<11161> A_IWL<11160> A_IWL<11159> A_IWL<11158> A_IWL<11157> A_IWL<11156> A_IWL<11155> A_IWL<11154> A_IWL<11153> A_IWL<11152> A_IWL<11151> A_IWL<11150> A_IWL<11149> A_IWL<11148> A_IWL<11147> A_IWL<11146> A_IWL<11145> A_IWL<11144> A_IWL<11143> A_IWL<11142> A_IWL<11141> A_IWL<11140> A_IWL<11139> A_IWL<11138> A_IWL<11137> A_IWL<11136> A_IWL<11135> A_IWL<11134> A_IWL<11133> A_IWL<11132> A_IWL<11131> A_IWL<11130> A_IWL<11129> A_IWL<11128> A_IWL<11127> A_IWL<11126> A_IWL<11125> A_IWL<11124> A_IWL<11123> A_IWL<11122> A_IWL<11121> A_IWL<11120> A_IWL<11119> A_IWL<11118> A_IWL<11117> A_IWL<11116> A_IWL<11115> A_IWL<11114> A_IWL<11113> A_IWL<11112> A_IWL<11111> A_IWL<11110> A_IWL<11109> A_IWL<11108> A_IWL<11107> A_IWL<11106> A_IWL<11105> A_IWL<11104> A_IWL<11103> A_IWL<11102> A_IWL<11101> A_IWL<11100> A_IWL<11099> A_IWL<11098> A_IWL<11097> A_IWL<11096> A_IWL<11095> A_IWL<11094> A_IWL<11093> A_IWL<11092> A_IWL<11091> A_IWL<11090> A_IWL<11089> A_IWL<11088> A_IWL<11087> A_IWL<11086> A_IWL<11085> A_IWL<11084> A_IWL<11083> A_IWL<11082> A_IWL<11081> A_IWL<11080> A_IWL<11079> A_IWL<11078> A_IWL<11077> A_IWL<11076> A_IWL<11075> A_IWL<11074> A_IWL<11073> A_IWL<11072> A_IWL<11071> A_IWL<11070> A_IWL<11069> A_IWL<11068> A_IWL<11067> A_IWL<11066> A_IWL<11065> A_IWL<11064> A_IWL<11063> A_IWL<11062> A_IWL<11061> A_IWL<11060> A_IWL<11059> A_IWL<11058> A_IWL<11057> A_IWL<11056> A_IWL<11055> A_IWL<11054> A_IWL<11053> A_IWL<11052> A_IWL<11051> A_IWL<11050> A_IWL<11049> A_IWL<11048> A_IWL<11047> A_IWL<11046> A_IWL<11045> A_IWL<11044> A_IWL<11043> A_IWL<11042> A_IWL<11041> A_IWL<11040> A_IWL<11039> A_IWL<11038> A_IWL<11037> A_IWL<11036> A_IWL<11035> A_IWL<11034> A_IWL<11033> A_IWL<11032> A_IWL<11031> A_IWL<11030> A_IWL<11029> A_IWL<11028> A_IWL<11027> A_IWL<11026> A_IWL<11025> A_IWL<11024> A_IWL<11023> A_IWL<11022> A_IWL<11021> A_IWL<11020> A_IWL<11019> A_IWL<11018> A_IWL<11017> A_IWL<11016> A_IWL<11015> A_IWL<11014> A_IWL<11013> A_IWL<11012> A_IWL<11011> A_IWL<11010> A_IWL<11009> A_IWL<11008> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<42> A_BLC<85> A_BLC<84> A_BLC_TOP<85> A_BLC_TOP<84> A_BLT<85> A_BLT<84> A_BLT_TOP<85> A_BLT_TOP<84> A_IWL<10751> A_IWL<10750> A_IWL<10749> A_IWL<10748> A_IWL<10747> A_IWL<10746> A_IWL<10745> A_IWL<10744> A_IWL<10743> A_IWL<10742> A_IWL<10741> A_IWL<10740> A_IWL<10739> A_IWL<10738> A_IWL<10737> A_IWL<10736> A_IWL<10735> A_IWL<10734> A_IWL<10733> A_IWL<10732> A_IWL<10731> A_IWL<10730> A_IWL<10729> A_IWL<10728> A_IWL<10727> A_IWL<10726> A_IWL<10725> A_IWL<10724> A_IWL<10723> A_IWL<10722> A_IWL<10721> A_IWL<10720> A_IWL<10719> A_IWL<10718> A_IWL<10717> A_IWL<10716> A_IWL<10715> A_IWL<10714> A_IWL<10713> A_IWL<10712> A_IWL<10711> A_IWL<10710> A_IWL<10709> A_IWL<10708> A_IWL<10707> A_IWL<10706> A_IWL<10705> A_IWL<10704> A_IWL<10703> A_IWL<10702> A_IWL<10701> A_IWL<10700> A_IWL<10699> A_IWL<10698> A_IWL<10697> A_IWL<10696> A_IWL<10695> A_IWL<10694> A_IWL<10693> A_IWL<10692> A_IWL<10691> A_IWL<10690> A_IWL<10689> A_IWL<10688> A_IWL<10687> A_IWL<10686> A_IWL<10685> A_IWL<10684> A_IWL<10683> A_IWL<10682> A_IWL<10681> A_IWL<10680> A_IWL<10679> A_IWL<10678> A_IWL<10677> A_IWL<10676> A_IWL<10675> A_IWL<10674> A_IWL<10673> A_IWL<10672> A_IWL<10671> A_IWL<10670> A_IWL<10669> A_IWL<10668> A_IWL<10667> A_IWL<10666> A_IWL<10665> A_IWL<10664> A_IWL<10663> A_IWL<10662> A_IWL<10661> A_IWL<10660> A_IWL<10659> A_IWL<10658> A_IWL<10657> A_IWL<10656> A_IWL<10655> A_IWL<10654> A_IWL<10653> A_IWL<10652> A_IWL<10651> A_IWL<10650> A_IWL<10649> A_IWL<10648> A_IWL<10647> A_IWL<10646> A_IWL<10645> A_IWL<10644> A_IWL<10643> A_IWL<10642> A_IWL<10641> A_IWL<10640> A_IWL<10639> A_IWL<10638> A_IWL<10637> A_IWL<10636> A_IWL<10635> A_IWL<10634> A_IWL<10633> A_IWL<10632> A_IWL<10631> A_IWL<10630> A_IWL<10629> A_IWL<10628> A_IWL<10627> A_IWL<10626> A_IWL<10625> A_IWL<10624> A_IWL<10623> A_IWL<10622> A_IWL<10621> A_IWL<10620> A_IWL<10619> A_IWL<10618> A_IWL<10617> A_IWL<10616> A_IWL<10615> A_IWL<10614> A_IWL<10613> A_IWL<10612> A_IWL<10611> A_IWL<10610> A_IWL<10609> A_IWL<10608> A_IWL<10607> A_IWL<10606> A_IWL<10605> A_IWL<10604> A_IWL<10603> A_IWL<10602> A_IWL<10601> A_IWL<10600> A_IWL<10599> A_IWL<10598> A_IWL<10597> A_IWL<10596> A_IWL<10595> A_IWL<10594> A_IWL<10593> A_IWL<10592> A_IWL<10591> A_IWL<10590> A_IWL<10589> A_IWL<10588> A_IWL<10587> A_IWL<10586> A_IWL<10585> A_IWL<10584> A_IWL<10583> A_IWL<10582> A_IWL<10581> A_IWL<10580> A_IWL<10579> A_IWL<10578> A_IWL<10577> A_IWL<10576> A_IWL<10575> A_IWL<10574> A_IWL<10573> A_IWL<10572> A_IWL<10571> A_IWL<10570> A_IWL<10569> A_IWL<10568> A_IWL<10567> A_IWL<10566> A_IWL<10565> A_IWL<10564> A_IWL<10563> A_IWL<10562> A_IWL<10561> A_IWL<10560> A_IWL<10559> A_IWL<10558> A_IWL<10557> A_IWL<10556> A_IWL<10555> A_IWL<10554> A_IWL<10553> A_IWL<10552> A_IWL<10551> A_IWL<10550> A_IWL<10549> A_IWL<10548> A_IWL<10547> A_IWL<10546> A_IWL<10545> A_IWL<10544> A_IWL<10543> A_IWL<10542> A_IWL<10541> A_IWL<10540> A_IWL<10539> A_IWL<10538> A_IWL<10537> A_IWL<10536> A_IWL<10535> A_IWL<10534> A_IWL<10533> A_IWL<10532> A_IWL<10531> A_IWL<10530> A_IWL<10529> A_IWL<10528> A_IWL<10527> A_IWL<10526> A_IWL<10525> A_IWL<10524> A_IWL<10523> A_IWL<10522> A_IWL<10521> A_IWL<10520> A_IWL<10519> A_IWL<10518> A_IWL<10517> A_IWL<10516> A_IWL<10515> A_IWL<10514> A_IWL<10513> A_IWL<10512> A_IWL<10511> A_IWL<10510> A_IWL<10509> A_IWL<10508> A_IWL<10507> A_IWL<10506> A_IWL<10505> A_IWL<10504> A_IWL<10503> A_IWL<10502> A_IWL<10501> A_IWL<10500> A_IWL<10499> A_IWL<10498> A_IWL<10497> A_IWL<10496> A_IWL<11007> A_IWL<11006> A_IWL<11005> A_IWL<11004> A_IWL<11003> A_IWL<11002> A_IWL<11001> A_IWL<11000> A_IWL<10999> A_IWL<10998> A_IWL<10997> A_IWL<10996> A_IWL<10995> A_IWL<10994> A_IWL<10993> A_IWL<10992> A_IWL<10991> A_IWL<10990> A_IWL<10989> A_IWL<10988> A_IWL<10987> A_IWL<10986> A_IWL<10985> A_IWL<10984> A_IWL<10983> A_IWL<10982> A_IWL<10981> A_IWL<10980> A_IWL<10979> A_IWL<10978> A_IWL<10977> A_IWL<10976> A_IWL<10975> A_IWL<10974> A_IWL<10973> A_IWL<10972> A_IWL<10971> A_IWL<10970> A_IWL<10969> A_IWL<10968> A_IWL<10967> A_IWL<10966> A_IWL<10965> A_IWL<10964> A_IWL<10963> A_IWL<10962> A_IWL<10961> A_IWL<10960> A_IWL<10959> A_IWL<10958> A_IWL<10957> A_IWL<10956> A_IWL<10955> A_IWL<10954> A_IWL<10953> A_IWL<10952> A_IWL<10951> A_IWL<10950> A_IWL<10949> A_IWL<10948> A_IWL<10947> A_IWL<10946> A_IWL<10945> A_IWL<10944> A_IWL<10943> A_IWL<10942> A_IWL<10941> A_IWL<10940> A_IWL<10939> A_IWL<10938> A_IWL<10937> A_IWL<10936> A_IWL<10935> A_IWL<10934> A_IWL<10933> A_IWL<10932> A_IWL<10931> A_IWL<10930> A_IWL<10929> A_IWL<10928> A_IWL<10927> A_IWL<10926> A_IWL<10925> A_IWL<10924> A_IWL<10923> A_IWL<10922> A_IWL<10921> A_IWL<10920> A_IWL<10919> A_IWL<10918> A_IWL<10917> A_IWL<10916> A_IWL<10915> A_IWL<10914> A_IWL<10913> A_IWL<10912> A_IWL<10911> A_IWL<10910> A_IWL<10909> A_IWL<10908> A_IWL<10907> A_IWL<10906> A_IWL<10905> A_IWL<10904> A_IWL<10903> A_IWL<10902> A_IWL<10901> A_IWL<10900> A_IWL<10899> A_IWL<10898> A_IWL<10897> A_IWL<10896> A_IWL<10895> A_IWL<10894> A_IWL<10893> A_IWL<10892> A_IWL<10891> A_IWL<10890> A_IWL<10889> A_IWL<10888> A_IWL<10887> A_IWL<10886> A_IWL<10885> A_IWL<10884> A_IWL<10883> A_IWL<10882> A_IWL<10881> A_IWL<10880> A_IWL<10879> A_IWL<10878> A_IWL<10877> A_IWL<10876> A_IWL<10875> A_IWL<10874> A_IWL<10873> A_IWL<10872> A_IWL<10871> A_IWL<10870> A_IWL<10869> A_IWL<10868> A_IWL<10867> A_IWL<10866> A_IWL<10865> A_IWL<10864> A_IWL<10863> A_IWL<10862> A_IWL<10861> A_IWL<10860> A_IWL<10859> A_IWL<10858> A_IWL<10857> A_IWL<10856> A_IWL<10855> A_IWL<10854> A_IWL<10853> A_IWL<10852> A_IWL<10851> A_IWL<10850> A_IWL<10849> A_IWL<10848> A_IWL<10847> A_IWL<10846> A_IWL<10845> A_IWL<10844> A_IWL<10843> A_IWL<10842> A_IWL<10841> A_IWL<10840> A_IWL<10839> A_IWL<10838> A_IWL<10837> A_IWL<10836> A_IWL<10835> A_IWL<10834> A_IWL<10833> A_IWL<10832> A_IWL<10831> A_IWL<10830> A_IWL<10829> A_IWL<10828> A_IWL<10827> A_IWL<10826> A_IWL<10825> A_IWL<10824> A_IWL<10823> A_IWL<10822> A_IWL<10821> A_IWL<10820> A_IWL<10819> A_IWL<10818> A_IWL<10817> A_IWL<10816> A_IWL<10815> A_IWL<10814> A_IWL<10813> A_IWL<10812> A_IWL<10811> A_IWL<10810> A_IWL<10809> A_IWL<10808> A_IWL<10807> A_IWL<10806> A_IWL<10805> A_IWL<10804> A_IWL<10803> A_IWL<10802> A_IWL<10801> A_IWL<10800> A_IWL<10799> A_IWL<10798> A_IWL<10797> A_IWL<10796> A_IWL<10795> A_IWL<10794> A_IWL<10793> A_IWL<10792> A_IWL<10791> A_IWL<10790> A_IWL<10789> A_IWL<10788> A_IWL<10787> A_IWL<10786> A_IWL<10785> A_IWL<10784> A_IWL<10783> A_IWL<10782> A_IWL<10781> A_IWL<10780> A_IWL<10779> A_IWL<10778> A_IWL<10777> A_IWL<10776> A_IWL<10775> A_IWL<10774> A_IWL<10773> A_IWL<10772> A_IWL<10771> A_IWL<10770> A_IWL<10769> A_IWL<10768> A_IWL<10767> A_IWL<10766> A_IWL<10765> A_IWL<10764> A_IWL<10763> A_IWL<10762> A_IWL<10761> A_IWL<10760> A_IWL<10759> A_IWL<10758> A_IWL<10757> A_IWL<10756> A_IWL<10755> A_IWL<10754> A_IWL<10753> A_IWL<10752> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<41> A_BLC<83> A_BLC<82> A_BLC_TOP<83> A_BLC_TOP<82> A_BLT<83> A_BLT<82> A_BLT_TOP<83> A_BLT_TOP<82> A_IWL<10495> A_IWL<10494> A_IWL<10493> A_IWL<10492> A_IWL<10491> A_IWL<10490> A_IWL<10489> A_IWL<10488> A_IWL<10487> A_IWL<10486> A_IWL<10485> A_IWL<10484> A_IWL<10483> A_IWL<10482> A_IWL<10481> A_IWL<10480> A_IWL<10479> A_IWL<10478> A_IWL<10477> A_IWL<10476> A_IWL<10475> A_IWL<10474> A_IWL<10473> A_IWL<10472> A_IWL<10471> A_IWL<10470> A_IWL<10469> A_IWL<10468> A_IWL<10467> A_IWL<10466> A_IWL<10465> A_IWL<10464> A_IWL<10463> A_IWL<10462> A_IWL<10461> A_IWL<10460> A_IWL<10459> A_IWL<10458> A_IWL<10457> A_IWL<10456> A_IWL<10455> A_IWL<10454> A_IWL<10453> A_IWL<10452> A_IWL<10451> A_IWL<10450> A_IWL<10449> A_IWL<10448> A_IWL<10447> A_IWL<10446> A_IWL<10445> A_IWL<10444> A_IWL<10443> A_IWL<10442> A_IWL<10441> A_IWL<10440> A_IWL<10439> A_IWL<10438> A_IWL<10437> A_IWL<10436> A_IWL<10435> A_IWL<10434> A_IWL<10433> A_IWL<10432> A_IWL<10431> A_IWL<10430> A_IWL<10429> A_IWL<10428> A_IWL<10427> A_IWL<10426> A_IWL<10425> A_IWL<10424> A_IWL<10423> A_IWL<10422> A_IWL<10421> A_IWL<10420> A_IWL<10419> A_IWL<10418> A_IWL<10417> A_IWL<10416> A_IWL<10415> A_IWL<10414> A_IWL<10413> A_IWL<10412> A_IWL<10411> A_IWL<10410> A_IWL<10409> A_IWL<10408> A_IWL<10407> A_IWL<10406> A_IWL<10405> A_IWL<10404> A_IWL<10403> A_IWL<10402> A_IWL<10401> A_IWL<10400> A_IWL<10399> A_IWL<10398> A_IWL<10397> A_IWL<10396> A_IWL<10395> A_IWL<10394> A_IWL<10393> A_IWL<10392> A_IWL<10391> A_IWL<10390> A_IWL<10389> A_IWL<10388> A_IWL<10387> A_IWL<10386> A_IWL<10385> A_IWL<10384> A_IWL<10383> A_IWL<10382> A_IWL<10381> A_IWL<10380> A_IWL<10379> A_IWL<10378> A_IWL<10377> A_IWL<10376> A_IWL<10375> A_IWL<10374> A_IWL<10373> A_IWL<10372> A_IWL<10371> A_IWL<10370> A_IWL<10369> A_IWL<10368> A_IWL<10367> A_IWL<10366> A_IWL<10365> A_IWL<10364> A_IWL<10363> A_IWL<10362> A_IWL<10361> A_IWL<10360> A_IWL<10359> A_IWL<10358> A_IWL<10357> A_IWL<10356> A_IWL<10355> A_IWL<10354> A_IWL<10353> A_IWL<10352> A_IWL<10351> A_IWL<10350> A_IWL<10349> A_IWL<10348> A_IWL<10347> A_IWL<10346> A_IWL<10345> A_IWL<10344> A_IWL<10343> A_IWL<10342> A_IWL<10341> A_IWL<10340> A_IWL<10339> A_IWL<10338> A_IWL<10337> A_IWL<10336> A_IWL<10335> A_IWL<10334> A_IWL<10333> A_IWL<10332> A_IWL<10331> A_IWL<10330> A_IWL<10329> A_IWL<10328> A_IWL<10327> A_IWL<10326> A_IWL<10325> A_IWL<10324> A_IWL<10323> A_IWL<10322> A_IWL<10321> A_IWL<10320> A_IWL<10319> A_IWL<10318> A_IWL<10317> A_IWL<10316> A_IWL<10315> A_IWL<10314> A_IWL<10313> A_IWL<10312> A_IWL<10311> A_IWL<10310> A_IWL<10309> A_IWL<10308> A_IWL<10307> A_IWL<10306> A_IWL<10305> A_IWL<10304> A_IWL<10303> A_IWL<10302> A_IWL<10301> A_IWL<10300> A_IWL<10299> A_IWL<10298> A_IWL<10297> A_IWL<10296> A_IWL<10295> A_IWL<10294> A_IWL<10293> A_IWL<10292> A_IWL<10291> A_IWL<10290> A_IWL<10289> A_IWL<10288> A_IWL<10287> A_IWL<10286> A_IWL<10285> A_IWL<10284> A_IWL<10283> A_IWL<10282> A_IWL<10281> A_IWL<10280> A_IWL<10279> A_IWL<10278> A_IWL<10277> A_IWL<10276> A_IWL<10275> A_IWL<10274> A_IWL<10273> A_IWL<10272> A_IWL<10271> A_IWL<10270> A_IWL<10269> A_IWL<10268> A_IWL<10267> A_IWL<10266> A_IWL<10265> A_IWL<10264> A_IWL<10263> A_IWL<10262> A_IWL<10261> A_IWL<10260> A_IWL<10259> A_IWL<10258> A_IWL<10257> A_IWL<10256> A_IWL<10255> A_IWL<10254> A_IWL<10253> A_IWL<10252> A_IWL<10251> A_IWL<10250> A_IWL<10249> A_IWL<10248> A_IWL<10247> A_IWL<10246> A_IWL<10245> A_IWL<10244> A_IWL<10243> A_IWL<10242> A_IWL<10241> A_IWL<10240> A_IWL<10751> A_IWL<10750> A_IWL<10749> A_IWL<10748> A_IWL<10747> A_IWL<10746> A_IWL<10745> A_IWL<10744> A_IWL<10743> A_IWL<10742> A_IWL<10741> A_IWL<10740> A_IWL<10739> A_IWL<10738> A_IWL<10737> A_IWL<10736> A_IWL<10735> A_IWL<10734> A_IWL<10733> A_IWL<10732> A_IWL<10731> A_IWL<10730> A_IWL<10729> A_IWL<10728> A_IWL<10727> A_IWL<10726> A_IWL<10725> A_IWL<10724> A_IWL<10723> A_IWL<10722> A_IWL<10721> A_IWL<10720> A_IWL<10719> A_IWL<10718> A_IWL<10717> A_IWL<10716> A_IWL<10715> A_IWL<10714> A_IWL<10713> A_IWL<10712> A_IWL<10711> A_IWL<10710> A_IWL<10709> A_IWL<10708> A_IWL<10707> A_IWL<10706> A_IWL<10705> A_IWL<10704> A_IWL<10703> A_IWL<10702> A_IWL<10701> A_IWL<10700> A_IWL<10699> A_IWL<10698> A_IWL<10697> A_IWL<10696> A_IWL<10695> A_IWL<10694> A_IWL<10693> A_IWL<10692> A_IWL<10691> A_IWL<10690> A_IWL<10689> A_IWL<10688> A_IWL<10687> A_IWL<10686> A_IWL<10685> A_IWL<10684> A_IWL<10683> A_IWL<10682> A_IWL<10681> A_IWL<10680> A_IWL<10679> A_IWL<10678> A_IWL<10677> A_IWL<10676> A_IWL<10675> A_IWL<10674> A_IWL<10673> A_IWL<10672> A_IWL<10671> A_IWL<10670> A_IWL<10669> A_IWL<10668> A_IWL<10667> A_IWL<10666> A_IWL<10665> A_IWL<10664> A_IWL<10663> A_IWL<10662> A_IWL<10661> A_IWL<10660> A_IWL<10659> A_IWL<10658> A_IWL<10657> A_IWL<10656> A_IWL<10655> A_IWL<10654> A_IWL<10653> A_IWL<10652> A_IWL<10651> A_IWL<10650> A_IWL<10649> A_IWL<10648> A_IWL<10647> A_IWL<10646> A_IWL<10645> A_IWL<10644> A_IWL<10643> A_IWL<10642> A_IWL<10641> A_IWL<10640> A_IWL<10639> A_IWL<10638> A_IWL<10637> A_IWL<10636> A_IWL<10635> A_IWL<10634> A_IWL<10633> A_IWL<10632> A_IWL<10631> A_IWL<10630> A_IWL<10629> A_IWL<10628> A_IWL<10627> A_IWL<10626> A_IWL<10625> A_IWL<10624> A_IWL<10623> A_IWL<10622> A_IWL<10621> A_IWL<10620> A_IWL<10619> A_IWL<10618> A_IWL<10617> A_IWL<10616> A_IWL<10615> A_IWL<10614> A_IWL<10613> A_IWL<10612> A_IWL<10611> A_IWL<10610> A_IWL<10609> A_IWL<10608> A_IWL<10607> A_IWL<10606> A_IWL<10605> A_IWL<10604> A_IWL<10603> A_IWL<10602> A_IWL<10601> A_IWL<10600> A_IWL<10599> A_IWL<10598> A_IWL<10597> A_IWL<10596> A_IWL<10595> A_IWL<10594> A_IWL<10593> A_IWL<10592> A_IWL<10591> A_IWL<10590> A_IWL<10589> A_IWL<10588> A_IWL<10587> A_IWL<10586> A_IWL<10585> A_IWL<10584> A_IWL<10583> A_IWL<10582> A_IWL<10581> A_IWL<10580> A_IWL<10579> A_IWL<10578> A_IWL<10577> A_IWL<10576> A_IWL<10575> A_IWL<10574> A_IWL<10573> A_IWL<10572> A_IWL<10571> A_IWL<10570> A_IWL<10569> A_IWL<10568> A_IWL<10567> A_IWL<10566> A_IWL<10565> A_IWL<10564> A_IWL<10563> A_IWL<10562> A_IWL<10561> A_IWL<10560> A_IWL<10559> A_IWL<10558> A_IWL<10557> A_IWL<10556> A_IWL<10555> A_IWL<10554> A_IWL<10553> A_IWL<10552> A_IWL<10551> A_IWL<10550> A_IWL<10549> A_IWL<10548> A_IWL<10547> A_IWL<10546> A_IWL<10545> A_IWL<10544> A_IWL<10543> A_IWL<10542> A_IWL<10541> A_IWL<10540> A_IWL<10539> A_IWL<10538> A_IWL<10537> A_IWL<10536> A_IWL<10535> A_IWL<10534> A_IWL<10533> A_IWL<10532> A_IWL<10531> A_IWL<10530> A_IWL<10529> A_IWL<10528> A_IWL<10527> A_IWL<10526> A_IWL<10525> A_IWL<10524> A_IWL<10523> A_IWL<10522> A_IWL<10521> A_IWL<10520> A_IWL<10519> A_IWL<10518> A_IWL<10517> A_IWL<10516> A_IWL<10515> A_IWL<10514> A_IWL<10513> A_IWL<10512> A_IWL<10511> A_IWL<10510> A_IWL<10509> A_IWL<10508> A_IWL<10507> A_IWL<10506> A_IWL<10505> A_IWL<10504> A_IWL<10503> A_IWL<10502> A_IWL<10501> A_IWL<10500> A_IWL<10499> A_IWL<10498> A_IWL<10497> A_IWL<10496> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<40> A_BLC<81> A_BLC<80> A_BLC_TOP<81> A_BLC_TOP<80> A_BLT<81> A_BLT<80> A_BLT_TOP<81> A_BLT_TOP<80> A_IWL<10239> A_IWL<10238> A_IWL<10237> A_IWL<10236> A_IWL<10235> A_IWL<10234> A_IWL<10233> A_IWL<10232> A_IWL<10231> A_IWL<10230> A_IWL<10229> A_IWL<10228> A_IWL<10227> A_IWL<10226> A_IWL<10225> A_IWL<10224> A_IWL<10223> A_IWL<10222> A_IWL<10221> A_IWL<10220> A_IWL<10219> A_IWL<10218> A_IWL<10217> A_IWL<10216> A_IWL<10215> A_IWL<10214> A_IWL<10213> A_IWL<10212> A_IWL<10211> A_IWL<10210> A_IWL<10209> A_IWL<10208> A_IWL<10207> A_IWL<10206> A_IWL<10205> A_IWL<10204> A_IWL<10203> A_IWL<10202> A_IWL<10201> A_IWL<10200> A_IWL<10199> A_IWL<10198> A_IWL<10197> A_IWL<10196> A_IWL<10195> A_IWL<10194> A_IWL<10193> A_IWL<10192> A_IWL<10191> A_IWL<10190> A_IWL<10189> A_IWL<10188> A_IWL<10187> A_IWL<10186> A_IWL<10185> A_IWL<10184> A_IWL<10183> A_IWL<10182> A_IWL<10181> A_IWL<10180> A_IWL<10179> A_IWL<10178> A_IWL<10177> A_IWL<10176> A_IWL<10175> A_IWL<10174> A_IWL<10173> A_IWL<10172> A_IWL<10171> A_IWL<10170> A_IWL<10169> A_IWL<10168> A_IWL<10167> A_IWL<10166> A_IWL<10165> A_IWL<10164> A_IWL<10163> A_IWL<10162> A_IWL<10161> A_IWL<10160> A_IWL<10159> A_IWL<10158> A_IWL<10157> A_IWL<10156> A_IWL<10155> A_IWL<10154> A_IWL<10153> A_IWL<10152> A_IWL<10151> A_IWL<10150> A_IWL<10149> A_IWL<10148> A_IWL<10147> A_IWL<10146> A_IWL<10145> A_IWL<10144> A_IWL<10143> A_IWL<10142> A_IWL<10141> A_IWL<10140> A_IWL<10139> A_IWL<10138> A_IWL<10137> A_IWL<10136> A_IWL<10135> A_IWL<10134> A_IWL<10133> A_IWL<10132> A_IWL<10131> A_IWL<10130> A_IWL<10129> A_IWL<10128> A_IWL<10127> A_IWL<10126> A_IWL<10125> A_IWL<10124> A_IWL<10123> A_IWL<10122> A_IWL<10121> A_IWL<10120> A_IWL<10119> A_IWL<10118> A_IWL<10117> A_IWL<10116> A_IWL<10115> A_IWL<10114> A_IWL<10113> A_IWL<10112> A_IWL<10111> A_IWL<10110> A_IWL<10109> A_IWL<10108> A_IWL<10107> A_IWL<10106> A_IWL<10105> A_IWL<10104> A_IWL<10103> A_IWL<10102> A_IWL<10101> A_IWL<10100> A_IWL<10099> A_IWL<10098> A_IWL<10097> A_IWL<10096> A_IWL<10095> A_IWL<10094> A_IWL<10093> A_IWL<10092> A_IWL<10091> A_IWL<10090> A_IWL<10089> A_IWL<10088> A_IWL<10087> A_IWL<10086> A_IWL<10085> A_IWL<10084> A_IWL<10083> A_IWL<10082> A_IWL<10081> A_IWL<10080> A_IWL<10079> A_IWL<10078> A_IWL<10077> A_IWL<10076> A_IWL<10075> A_IWL<10074> A_IWL<10073> A_IWL<10072> A_IWL<10071> A_IWL<10070> A_IWL<10069> A_IWL<10068> A_IWL<10067> A_IWL<10066> A_IWL<10065> A_IWL<10064> A_IWL<10063> A_IWL<10062> A_IWL<10061> A_IWL<10060> A_IWL<10059> A_IWL<10058> A_IWL<10057> A_IWL<10056> A_IWL<10055> A_IWL<10054> A_IWL<10053> A_IWL<10052> A_IWL<10051> A_IWL<10050> A_IWL<10049> A_IWL<10048> A_IWL<10047> A_IWL<10046> A_IWL<10045> A_IWL<10044> A_IWL<10043> A_IWL<10042> A_IWL<10041> A_IWL<10040> A_IWL<10039> A_IWL<10038> A_IWL<10037> A_IWL<10036> A_IWL<10035> A_IWL<10034> A_IWL<10033> A_IWL<10032> A_IWL<10031> A_IWL<10030> A_IWL<10029> A_IWL<10028> A_IWL<10027> A_IWL<10026> A_IWL<10025> A_IWL<10024> A_IWL<10023> A_IWL<10022> A_IWL<10021> A_IWL<10020> A_IWL<10019> A_IWL<10018> A_IWL<10017> A_IWL<10016> A_IWL<10015> A_IWL<10014> A_IWL<10013> A_IWL<10012> A_IWL<10011> A_IWL<10010> A_IWL<10009> A_IWL<10008> A_IWL<10007> A_IWL<10006> A_IWL<10005> A_IWL<10004> A_IWL<10003> A_IWL<10002> A_IWL<10001> A_IWL<10000> A_IWL<9999> A_IWL<9998> A_IWL<9997> A_IWL<9996> A_IWL<9995> A_IWL<9994> A_IWL<9993> A_IWL<9992> A_IWL<9991> A_IWL<9990> A_IWL<9989> A_IWL<9988> A_IWL<9987> A_IWL<9986> A_IWL<9985> A_IWL<9984> A_IWL<10495> A_IWL<10494> A_IWL<10493> A_IWL<10492> A_IWL<10491> A_IWL<10490> A_IWL<10489> A_IWL<10488> A_IWL<10487> A_IWL<10486> A_IWL<10485> A_IWL<10484> A_IWL<10483> A_IWL<10482> A_IWL<10481> A_IWL<10480> A_IWL<10479> A_IWL<10478> A_IWL<10477> A_IWL<10476> A_IWL<10475> A_IWL<10474> A_IWL<10473> A_IWL<10472> A_IWL<10471> A_IWL<10470> A_IWL<10469> A_IWL<10468> A_IWL<10467> A_IWL<10466> A_IWL<10465> A_IWL<10464> A_IWL<10463> A_IWL<10462> A_IWL<10461> A_IWL<10460> A_IWL<10459> A_IWL<10458> A_IWL<10457> A_IWL<10456> A_IWL<10455> A_IWL<10454> A_IWL<10453> A_IWL<10452> A_IWL<10451> A_IWL<10450> A_IWL<10449> A_IWL<10448> A_IWL<10447> A_IWL<10446> A_IWL<10445> A_IWL<10444> A_IWL<10443> A_IWL<10442> A_IWL<10441> A_IWL<10440> A_IWL<10439> A_IWL<10438> A_IWL<10437> A_IWL<10436> A_IWL<10435> A_IWL<10434> A_IWL<10433> A_IWL<10432> A_IWL<10431> A_IWL<10430> A_IWL<10429> A_IWL<10428> A_IWL<10427> A_IWL<10426> A_IWL<10425> A_IWL<10424> A_IWL<10423> A_IWL<10422> A_IWL<10421> A_IWL<10420> A_IWL<10419> A_IWL<10418> A_IWL<10417> A_IWL<10416> A_IWL<10415> A_IWL<10414> A_IWL<10413> A_IWL<10412> A_IWL<10411> A_IWL<10410> A_IWL<10409> A_IWL<10408> A_IWL<10407> A_IWL<10406> A_IWL<10405> A_IWL<10404> A_IWL<10403> A_IWL<10402> A_IWL<10401> A_IWL<10400> A_IWL<10399> A_IWL<10398> A_IWL<10397> A_IWL<10396> A_IWL<10395> A_IWL<10394> A_IWL<10393> A_IWL<10392> A_IWL<10391> A_IWL<10390> A_IWL<10389> A_IWL<10388> A_IWL<10387> A_IWL<10386> A_IWL<10385> A_IWL<10384> A_IWL<10383> A_IWL<10382> A_IWL<10381> A_IWL<10380> A_IWL<10379> A_IWL<10378> A_IWL<10377> A_IWL<10376> A_IWL<10375> A_IWL<10374> A_IWL<10373> A_IWL<10372> A_IWL<10371> A_IWL<10370> A_IWL<10369> A_IWL<10368> A_IWL<10367> A_IWL<10366> A_IWL<10365> A_IWL<10364> A_IWL<10363> A_IWL<10362> A_IWL<10361> A_IWL<10360> A_IWL<10359> A_IWL<10358> A_IWL<10357> A_IWL<10356> A_IWL<10355> A_IWL<10354> A_IWL<10353> A_IWL<10352> A_IWL<10351> A_IWL<10350> A_IWL<10349> A_IWL<10348> A_IWL<10347> A_IWL<10346> A_IWL<10345> A_IWL<10344> A_IWL<10343> A_IWL<10342> A_IWL<10341> A_IWL<10340> A_IWL<10339> A_IWL<10338> A_IWL<10337> A_IWL<10336> A_IWL<10335> A_IWL<10334> A_IWL<10333> A_IWL<10332> A_IWL<10331> A_IWL<10330> A_IWL<10329> A_IWL<10328> A_IWL<10327> A_IWL<10326> A_IWL<10325> A_IWL<10324> A_IWL<10323> A_IWL<10322> A_IWL<10321> A_IWL<10320> A_IWL<10319> A_IWL<10318> A_IWL<10317> A_IWL<10316> A_IWL<10315> A_IWL<10314> A_IWL<10313> A_IWL<10312> A_IWL<10311> A_IWL<10310> A_IWL<10309> A_IWL<10308> A_IWL<10307> A_IWL<10306> A_IWL<10305> A_IWL<10304> A_IWL<10303> A_IWL<10302> A_IWL<10301> A_IWL<10300> A_IWL<10299> A_IWL<10298> A_IWL<10297> A_IWL<10296> A_IWL<10295> A_IWL<10294> A_IWL<10293> A_IWL<10292> A_IWL<10291> A_IWL<10290> A_IWL<10289> A_IWL<10288> A_IWL<10287> A_IWL<10286> A_IWL<10285> A_IWL<10284> A_IWL<10283> A_IWL<10282> A_IWL<10281> A_IWL<10280> A_IWL<10279> A_IWL<10278> A_IWL<10277> A_IWL<10276> A_IWL<10275> A_IWL<10274> A_IWL<10273> A_IWL<10272> A_IWL<10271> A_IWL<10270> A_IWL<10269> A_IWL<10268> A_IWL<10267> A_IWL<10266> A_IWL<10265> A_IWL<10264> A_IWL<10263> A_IWL<10262> A_IWL<10261> A_IWL<10260> A_IWL<10259> A_IWL<10258> A_IWL<10257> A_IWL<10256> A_IWL<10255> A_IWL<10254> A_IWL<10253> A_IWL<10252> A_IWL<10251> A_IWL<10250> A_IWL<10249> A_IWL<10248> A_IWL<10247> A_IWL<10246> A_IWL<10245> A_IWL<10244> A_IWL<10243> A_IWL<10242> A_IWL<10241> A_IWL<10240> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<39> A_BLC<79> A_BLC<78> A_BLC_TOP<79> A_BLC_TOP<78> A_BLT<79> A_BLT<78> A_BLT_TOP<79> A_BLT_TOP<78> A_IWL<9983> A_IWL<9982> A_IWL<9981> A_IWL<9980> A_IWL<9979> A_IWL<9978> A_IWL<9977> A_IWL<9976> A_IWL<9975> A_IWL<9974> A_IWL<9973> A_IWL<9972> A_IWL<9971> A_IWL<9970> A_IWL<9969> A_IWL<9968> A_IWL<9967> A_IWL<9966> A_IWL<9965> A_IWL<9964> A_IWL<9963> A_IWL<9962> A_IWL<9961> A_IWL<9960> A_IWL<9959> A_IWL<9958> A_IWL<9957> A_IWL<9956> A_IWL<9955> A_IWL<9954> A_IWL<9953> A_IWL<9952> A_IWL<9951> A_IWL<9950> A_IWL<9949> A_IWL<9948> A_IWL<9947> A_IWL<9946> A_IWL<9945> A_IWL<9944> A_IWL<9943> A_IWL<9942> A_IWL<9941> A_IWL<9940> A_IWL<9939> A_IWL<9938> A_IWL<9937> A_IWL<9936> A_IWL<9935> A_IWL<9934> A_IWL<9933> A_IWL<9932> A_IWL<9931> A_IWL<9930> A_IWL<9929> A_IWL<9928> A_IWL<9927> A_IWL<9926> A_IWL<9925> A_IWL<9924> A_IWL<9923> A_IWL<9922> A_IWL<9921> A_IWL<9920> A_IWL<9919> A_IWL<9918> A_IWL<9917> A_IWL<9916> A_IWL<9915> A_IWL<9914> A_IWL<9913> A_IWL<9912> A_IWL<9911> A_IWL<9910> A_IWL<9909> A_IWL<9908> A_IWL<9907> A_IWL<9906> A_IWL<9905> A_IWL<9904> A_IWL<9903> A_IWL<9902> A_IWL<9901> A_IWL<9900> A_IWL<9899> A_IWL<9898> A_IWL<9897> A_IWL<9896> A_IWL<9895> A_IWL<9894> A_IWL<9893> A_IWL<9892> A_IWL<9891> A_IWL<9890> A_IWL<9889> A_IWL<9888> A_IWL<9887> A_IWL<9886> A_IWL<9885> A_IWL<9884> A_IWL<9883> A_IWL<9882> A_IWL<9881> A_IWL<9880> A_IWL<9879> A_IWL<9878> A_IWL<9877> A_IWL<9876> A_IWL<9875> A_IWL<9874> A_IWL<9873> A_IWL<9872> A_IWL<9871> A_IWL<9870> A_IWL<9869> A_IWL<9868> A_IWL<9867> A_IWL<9866> A_IWL<9865> A_IWL<9864> A_IWL<9863> A_IWL<9862> A_IWL<9861> A_IWL<9860> A_IWL<9859> A_IWL<9858> A_IWL<9857> A_IWL<9856> A_IWL<9855> A_IWL<9854> A_IWL<9853> A_IWL<9852> A_IWL<9851> A_IWL<9850> A_IWL<9849> A_IWL<9848> A_IWL<9847> A_IWL<9846> A_IWL<9845> A_IWL<9844> A_IWL<9843> A_IWL<9842> A_IWL<9841> A_IWL<9840> A_IWL<9839> A_IWL<9838> A_IWL<9837> A_IWL<9836> A_IWL<9835> A_IWL<9834> A_IWL<9833> A_IWL<9832> A_IWL<9831> A_IWL<9830> A_IWL<9829> A_IWL<9828> A_IWL<9827> A_IWL<9826> A_IWL<9825> A_IWL<9824> A_IWL<9823> A_IWL<9822> A_IWL<9821> A_IWL<9820> A_IWL<9819> A_IWL<9818> A_IWL<9817> A_IWL<9816> A_IWL<9815> A_IWL<9814> A_IWL<9813> A_IWL<9812> A_IWL<9811> A_IWL<9810> A_IWL<9809> A_IWL<9808> A_IWL<9807> A_IWL<9806> A_IWL<9805> A_IWL<9804> A_IWL<9803> A_IWL<9802> A_IWL<9801> A_IWL<9800> A_IWL<9799> A_IWL<9798> A_IWL<9797> A_IWL<9796> A_IWL<9795> A_IWL<9794> A_IWL<9793> A_IWL<9792> A_IWL<9791> A_IWL<9790> A_IWL<9789> A_IWL<9788> A_IWL<9787> A_IWL<9786> A_IWL<9785> A_IWL<9784> A_IWL<9783> A_IWL<9782> A_IWL<9781> A_IWL<9780> A_IWL<9779> A_IWL<9778> A_IWL<9777> A_IWL<9776> A_IWL<9775> A_IWL<9774> A_IWL<9773> A_IWL<9772> A_IWL<9771> A_IWL<9770> A_IWL<9769> A_IWL<9768> A_IWL<9767> A_IWL<9766> A_IWL<9765> A_IWL<9764> A_IWL<9763> A_IWL<9762> A_IWL<9761> A_IWL<9760> A_IWL<9759> A_IWL<9758> A_IWL<9757> A_IWL<9756> A_IWL<9755> A_IWL<9754> A_IWL<9753> A_IWL<9752> A_IWL<9751> A_IWL<9750> A_IWL<9749> A_IWL<9748> A_IWL<9747> A_IWL<9746> A_IWL<9745> A_IWL<9744> A_IWL<9743> A_IWL<9742> A_IWL<9741> A_IWL<9740> A_IWL<9739> A_IWL<9738> A_IWL<9737> A_IWL<9736> A_IWL<9735> A_IWL<9734> A_IWL<9733> A_IWL<9732> A_IWL<9731> A_IWL<9730> A_IWL<9729> A_IWL<9728> A_IWL<10239> A_IWL<10238> A_IWL<10237> A_IWL<10236> A_IWL<10235> A_IWL<10234> A_IWL<10233> A_IWL<10232> A_IWL<10231> A_IWL<10230> A_IWL<10229> A_IWL<10228> A_IWL<10227> A_IWL<10226> A_IWL<10225> A_IWL<10224> A_IWL<10223> A_IWL<10222> A_IWL<10221> A_IWL<10220> A_IWL<10219> A_IWL<10218> A_IWL<10217> A_IWL<10216> A_IWL<10215> A_IWL<10214> A_IWL<10213> A_IWL<10212> A_IWL<10211> A_IWL<10210> A_IWL<10209> A_IWL<10208> A_IWL<10207> A_IWL<10206> A_IWL<10205> A_IWL<10204> A_IWL<10203> A_IWL<10202> A_IWL<10201> A_IWL<10200> A_IWL<10199> A_IWL<10198> A_IWL<10197> A_IWL<10196> A_IWL<10195> A_IWL<10194> A_IWL<10193> A_IWL<10192> A_IWL<10191> A_IWL<10190> A_IWL<10189> A_IWL<10188> A_IWL<10187> A_IWL<10186> A_IWL<10185> A_IWL<10184> A_IWL<10183> A_IWL<10182> A_IWL<10181> A_IWL<10180> A_IWL<10179> A_IWL<10178> A_IWL<10177> A_IWL<10176> A_IWL<10175> A_IWL<10174> A_IWL<10173> A_IWL<10172> A_IWL<10171> A_IWL<10170> A_IWL<10169> A_IWL<10168> A_IWL<10167> A_IWL<10166> A_IWL<10165> A_IWL<10164> A_IWL<10163> A_IWL<10162> A_IWL<10161> A_IWL<10160> A_IWL<10159> A_IWL<10158> A_IWL<10157> A_IWL<10156> A_IWL<10155> A_IWL<10154> A_IWL<10153> A_IWL<10152> A_IWL<10151> A_IWL<10150> A_IWL<10149> A_IWL<10148> A_IWL<10147> A_IWL<10146> A_IWL<10145> A_IWL<10144> A_IWL<10143> A_IWL<10142> A_IWL<10141> A_IWL<10140> A_IWL<10139> A_IWL<10138> A_IWL<10137> A_IWL<10136> A_IWL<10135> A_IWL<10134> A_IWL<10133> A_IWL<10132> A_IWL<10131> A_IWL<10130> A_IWL<10129> A_IWL<10128> A_IWL<10127> A_IWL<10126> A_IWL<10125> A_IWL<10124> A_IWL<10123> A_IWL<10122> A_IWL<10121> A_IWL<10120> A_IWL<10119> A_IWL<10118> A_IWL<10117> A_IWL<10116> A_IWL<10115> A_IWL<10114> A_IWL<10113> A_IWL<10112> A_IWL<10111> A_IWL<10110> A_IWL<10109> A_IWL<10108> A_IWL<10107> A_IWL<10106> A_IWL<10105> A_IWL<10104> A_IWL<10103> A_IWL<10102> A_IWL<10101> A_IWL<10100> A_IWL<10099> A_IWL<10098> A_IWL<10097> A_IWL<10096> A_IWL<10095> A_IWL<10094> A_IWL<10093> A_IWL<10092> A_IWL<10091> A_IWL<10090> A_IWL<10089> A_IWL<10088> A_IWL<10087> A_IWL<10086> A_IWL<10085> A_IWL<10084> A_IWL<10083> A_IWL<10082> A_IWL<10081> A_IWL<10080> A_IWL<10079> A_IWL<10078> A_IWL<10077> A_IWL<10076> A_IWL<10075> A_IWL<10074> A_IWL<10073> A_IWL<10072> A_IWL<10071> A_IWL<10070> A_IWL<10069> A_IWL<10068> A_IWL<10067> A_IWL<10066> A_IWL<10065> A_IWL<10064> A_IWL<10063> A_IWL<10062> A_IWL<10061> A_IWL<10060> A_IWL<10059> A_IWL<10058> A_IWL<10057> A_IWL<10056> A_IWL<10055> A_IWL<10054> A_IWL<10053> A_IWL<10052> A_IWL<10051> A_IWL<10050> A_IWL<10049> A_IWL<10048> A_IWL<10047> A_IWL<10046> A_IWL<10045> A_IWL<10044> A_IWL<10043> A_IWL<10042> A_IWL<10041> A_IWL<10040> A_IWL<10039> A_IWL<10038> A_IWL<10037> A_IWL<10036> A_IWL<10035> A_IWL<10034> A_IWL<10033> A_IWL<10032> A_IWL<10031> A_IWL<10030> A_IWL<10029> A_IWL<10028> A_IWL<10027> A_IWL<10026> A_IWL<10025> A_IWL<10024> A_IWL<10023> A_IWL<10022> A_IWL<10021> A_IWL<10020> A_IWL<10019> A_IWL<10018> A_IWL<10017> A_IWL<10016> A_IWL<10015> A_IWL<10014> A_IWL<10013> A_IWL<10012> A_IWL<10011> A_IWL<10010> A_IWL<10009> A_IWL<10008> A_IWL<10007> A_IWL<10006> A_IWL<10005> A_IWL<10004> A_IWL<10003> A_IWL<10002> A_IWL<10001> A_IWL<10000> A_IWL<9999> A_IWL<9998> A_IWL<9997> A_IWL<9996> A_IWL<9995> A_IWL<9994> A_IWL<9993> A_IWL<9992> A_IWL<9991> A_IWL<9990> A_IWL<9989> A_IWL<9988> A_IWL<9987> A_IWL<9986> A_IWL<9985> A_IWL<9984> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<38> A_BLC<77> A_BLC<76> A_BLC_TOP<77> A_BLC_TOP<76> A_BLT<77> A_BLT<76> A_BLT_TOP<77> A_BLT_TOP<76> A_IWL<9727> A_IWL<9726> A_IWL<9725> A_IWL<9724> A_IWL<9723> A_IWL<9722> A_IWL<9721> A_IWL<9720> A_IWL<9719> A_IWL<9718> A_IWL<9717> A_IWL<9716> A_IWL<9715> A_IWL<9714> A_IWL<9713> A_IWL<9712> A_IWL<9711> A_IWL<9710> A_IWL<9709> A_IWL<9708> A_IWL<9707> A_IWL<9706> A_IWL<9705> A_IWL<9704> A_IWL<9703> A_IWL<9702> A_IWL<9701> A_IWL<9700> A_IWL<9699> A_IWL<9698> A_IWL<9697> A_IWL<9696> A_IWL<9695> A_IWL<9694> A_IWL<9693> A_IWL<9692> A_IWL<9691> A_IWL<9690> A_IWL<9689> A_IWL<9688> A_IWL<9687> A_IWL<9686> A_IWL<9685> A_IWL<9684> A_IWL<9683> A_IWL<9682> A_IWL<9681> A_IWL<9680> A_IWL<9679> A_IWL<9678> A_IWL<9677> A_IWL<9676> A_IWL<9675> A_IWL<9674> A_IWL<9673> A_IWL<9672> A_IWL<9671> A_IWL<9670> A_IWL<9669> A_IWL<9668> A_IWL<9667> A_IWL<9666> A_IWL<9665> A_IWL<9664> A_IWL<9663> A_IWL<9662> A_IWL<9661> A_IWL<9660> A_IWL<9659> A_IWL<9658> A_IWL<9657> A_IWL<9656> A_IWL<9655> A_IWL<9654> A_IWL<9653> A_IWL<9652> A_IWL<9651> A_IWL<9650> A_IWL<9649> A_IWL<9648> A_IWL<9647> A_IWL<9646> A_IWL<9645> A_IWL<9644> A_IWL<9643> A_IWL<9642> A_IWL<9641> A_IWL<9640> A_IWL<9639> A_IWL<9638> A_IWL<9637> A_IWL<9636> A_IWL<9635> A_IWL<9634> A_IWL<9633> A_IWL<9632> A_IWL<9631> A_IWL<9630> A_IWL<9629> A_IWL<9628> A_IWL<9627> A_IWL<9626> A_IWL<9625> A_IWL<9624> A_IWL<9623> A_IWL<9622> A_IWL<9621> A_IWL<9620> A_IWL<9619> A_IWL<9618> A_IWL<9617> A_IWL<9616> A_IWL<9615> A_IWL<9614> A_IWL<9613> A_IWL<9612> A_IWL<9611> A_IWL<9610> A_IWL<9609> A_IWL<9608> A_IWL<9607> A_IWL<9606> A_IWL<9605> A_IWL<9604> A_IWL<9603> A_IWL<9602> A_IWL<9601> A_IWL<9600> A_IWL<9599> A_IWL<9598> A_IWL<9597> A_IWL<9596> A_IWL<9595> A_IWL<9594> A_IWL<9593> A_IWL<9592> A_IWL<9591> A_IWL<9590> A_IWL<9589> A_IWL<9588> A_IWL<9587> A_IWL<9586> A_IWL<9585> A_IWL<9584> A_IWL<9583> A_IWL<9582> A_IWL<9581> A_IWL<9580> A_IWL<9579> A_IWL<9578> A_IWL<9577> A_IWL<9576> A_IWL<9575> A_IWL<9574> A_IWL<9573> A_IWL<9572> A_IWL<9571> A_IWL<9570> A_IWL<9569> A_IWL<9568> A_IWL<9567> A_IWL<9566> A_IWL<9565> A_IWL<9564> A_IWL<9563> A_IWL<9562> A_IWL<9561> A_IWL<9560> A_IWL<9559> A_IWL<9558> A_IWL<9557> A_IWL<9556> A_IWL<9555> A_IWL<9554> A_IWL<9553> A_IWL<9552> A_IWL<9551> A_IWL<9550> A_IWL<9549> A_IWL<9548> A_IWL<9547> A_IWL<9546> A_IWL<9545> A_IWL<9544> A_IWL<9543> A_IWL<9542> A_IWL<9541> A_IWL<9540> A_IWL<9539> A_IWL<9538> A_IWL<9537> A_IWL<9536> A_IWL<9535> A_IWL<9534> A_IWL<9533> A_IWL<9532> A_IWL<9531> A_IWL<9530> A_IWL<9529> A_IWL<9528> A_IWL<9527> A_IWL<9526> A_IWL<9525> A_IWL<9524> A_IWL<9523> A_IWL<9522> A_IWL<9521> A_IWL<9520> A_IWL<9519> A_IWL<9518> A_IWL<9517> A_IWL<9516> A_IWL<9515> A_IWL<9514> A_IWL<9513> A_IWL<9512> A_IWL<9511> A_IWL<9510> A_IWL<9509> A_IWL<9508> A_IWL<9507> A_IWL<9506> A_IWL<9505> A_IWL<9504> A_IWL<9503> A_IWL<9502> A_IWL<9501> A_IWL<9500> A_IWL<9499> A_IWL<9498> A_IWL<9497> A_IWL<9496> A_IWL<9495> A_IWL<9494> A_IWL<9493> A_IWL<9492> A_IWL<9491> A_IWL<9490> A_IWL<9489> A_IWL<9488> A_IWL<9487> A_IWL<9486> A_IWL<9485> A_IWL<9484> A_IWL<9483> A_IWL<9482> A_IWL<9481> A_IWL<9480> A_IWL<9479> A_IWL<9478> A_IWL<9477> A_IWL<9476> A_IWL<9475> A_IWL<9474> A_IWL<9473> A_IWL<9472> A_IWL<9983> A_IWL<9982> A_IWL<9981> A_IWL<9980> A_IWL<9979> A_IWL<9978> A_IWL<9977> A_IWL<9976> A_IWL<9975> A_IWL<9974> A_IWL<9973> A_IWL<9972> A_IWL<9971> A_IWL<9970> A_IWL<9969> A_IWL<9968> A_IWL<9967> A_IWL<9966> A_IWL<9965> A_IWL<9964> A_IWL<9963> A_IWL<9962> A_IWL<9961> A_IWL<9960> A_IWL<9959> A_IWL<9958> A_IWL<9957> A_IWL<9956> A_IWL<9955> A_IWL<9954> A_IWL<9953> A_IWL<9952> A_IWL<9951> A_IWL<9950> A_IWL<9949> A_IWL<9948> A_IWL<9947> A_IWL<9946> A_IWL<9945> A_IWL<9944> A_IWL<9943> A_IWL<9942> A_IWL<9941> A_IWL<9940> A_IWL<9939> A_IWL<9938> A_IWL<9937> A_IWL<9936> A_IWL<9935> A_IWL<9934> A_IWL<9933> A_IWL<9932> A_IWL<9931> A_IWL<9930> A_IWL<9929> A_IWL<9928> A_IWL<9927> A_IWL<9926> A_IWL<9925> A_IWL<9924> A_IWL<9923> A_IWL<9922> A_IWL<9921> A_IWL<9920> A_IWL<9919> A_IWL<9918> A_IWL<9917> A_IWL<9916> A_IWL<9915> A_IWL<9914> A_IWL<9913> A_IWL<9912> A_IWL<9911> A_IWL<9910> A_IWL<9909> A_IWL<9908> A_IWL<9907> A_IWL<9906> A_IWL<9905> A_IWL<9904> A_IWL<9903> A_IWL<9902> A_IWL<9901> A_IWL<9900> A_IWL<9899> A_IWL<9898> A_IWL<9897> A_IWL<9896> A_IWL<9895> A_IWL<9894> A_IWL<9893> A_IWL<9892> A_IWL<9891> A_IWL<9890> A_IWL<9889> A_IWL<9888> A_IWL<9887> A_IWL<9886> A_IWL<9885> A_IWL<9884> A_IWL<9883> A_IWL<9882> A_IWL<9881> A_IWL<9880> A_IWL<9879> A_IWL<9878> A_IWL<9877> A_IWL<9876> A_IWL<9875> A_IWL<9874> A_IWL<9873> A_IWL<9872> A_IWL<9871> A_IWL<9870> A_IWL<9869> A_IWL<9868> A_IWL<9867> A_IWL<9866> A_IWL<9865> A_IWL<9864> A_IWL<9863> A_IWL<9862> A_IWL<9861> A_IWL<9860> A_IWL<9859> A_IWL<9858> A_IWL<9857> A_IWL<9856> A_IWL<9855> A_IWL<9854> A_IWL<9853> A_IWL<9852> A_IWL<9851> A_IWL<9850> A_IWL<9849> A_IWL<9848> A_IWL<9847> A_IWL<9846> A_IWL<9845> A_IWL<9844> A_IWL<9843> A_IWL<9842> A_IWL<9841> A_IWL<9840> A_IWL<9839> A_IWL<9838> A_IWL<9837> A_IWL<9836> A_IWL<9835> A_IWL<9834> A_IWL<9833> A_IWL<9832> A_IWL<9831> A_IWL<9830> A_IWL<9829> A_IWL<9828> A_IWL<9827> A_IWL<9826> A_IWL<9825> A_IWL<9824> A_IWL<9823> A_IWL<9822> A_IWL<9821> A_IWL<9820> A_IWL<9819> A_IWL<9818> A_IWL<9817> A_IWL<9816> A_IWL<9815> A_IWL<9814> A_IWL<9813> A_IWL<9812> A_IWL<9811> A_IWL<9810> A_IWL<9809> A_IWL<9808> A_IWL<9807> A_IWL<9806> A_IWL<9805> A_IWL<9804> A_IWL<9803> A_IWL<9802> A_IWL<9801> A_IWL<9800> A_IWL<9799> A_IWL<9798> A_IWL<9797> A_IWL<9796> A_IWL<9795> A_IWL<9794> A_IWL<9793> A_IWL<9792> A_IWL<9791> A_IWL<9790> A_IWL<9789> A_IWL<9788> A_IWL<9787> A_IWL<9786> A_IWL<9785> A_IWL<9784> A_IWL<9783> A_IWL<9782> A_IWL<9781> A_IWL<9780> A_IWL<9779> A_IWL<9778> A_IWL<9777> A_IWL<9776> A_IWL<9775> A_IWL<9774> A_IWL<9773> A_IWL<9772> A_IWL<9771> A_IWL<9770> A_IWL<9769> A_IWL<9768> A_IWL<9767> A_IWL<9766> A_IWL<9765> A_IWL<9764> A_IWL<9763> A_IWL<9762> A_IWL<9761> A_IWL<9760> A_IWL<9759> A_IWL<9758> A_IWL<9757> A_IWL<9756> A_IWL<9755> A_IWL<9754> A_IWL<9753> A_IWL<9752> A_IWL<9751> A_IWL<9750> A_IWL<9749> A_IWL<9748> A_IWL<9747> A_IWL<9746> A_IWL<9745> A_IWL<9744> A_IWL<9743> A_IWL<9742> A_IWL<9741> A_IWL<9740> A_IWL<9739> A_IWL<9738> A_IWL<9737> A_IWL<9736> A_IWL<9735> A_IWL<9734> A_IWL<9733> A_IWL<9732> A_IWL<9731> A_IWL<9730> A_IWL<9729> A_IWL<9728> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<37> A_BLC<75> A_BLC<74> A_BLC_TOP<75> A_BLC_TOP<74> A_BLT<75> A_BLT<74> A_BLT_TOP<75> A_BLT_TOP<74> A_IWL<9471> A_IWL<9470> A_IWL<9469> A_IWL<9468> A_IWL<9467> A_IWL<9466> A_IWL<9465> A_IWL<9464> A_IWL<9463> A_IWL<9462> A_IWL<9461> A_IWL<9460> A_IWL<9459> A_IWL<9458> A_IWL<9457> A_IWL<9456> A_IWL<9455> A_IWL<9454> A_IWL<9453> A_IWL<9452> A_IWL<9451> A_IWL<9450> A_IWL<9449> A_IWL<9448> A_IWL<9447> A_IWL<9446> A_IWL<9445> A_IWL<9444> A_IWL<9443> A_IWL<9442> A_IWL<9441> A_IWL<9440> A_IWL<9439> A_IWL<9438> A_IWL<9437> A_IWL<9436> A_IWL<9435> A_IWL<9434> A_IWL<9433> A_IWL<9432> A_IWL<9431> A_IWL<9430> A_IWL<9429> A_IWL<9428> A_IWL<9427> A_IWL<9426> A_IWL<9425> A_IWL<9424> A_IWL<9423> A_IWL<9422> A_IWL<9421> A_IWL<9420> A_IWL<9419> A_IWL<9418> A_IWL<9417> A_IWL<9416> A_IWL<9415> A_IWL<9414> A_IWL<9413> A_IWL<9412> A_IWL<9411> A_IWL<9410> A_IWL<9409> A_IWL<9408> A_IWL<9407> A_IWL<9406> A_IWL<9405> A_IWL<9404> A_IWL<9403> A_IWL<9402> A_IWL<9401> A_IWL<9400> A_IWL<9399> A_IWL<9398> A_IWL<9397> A_IWL<9396> A_IWL<9395> A_IWL<9394> A_IWL<9393> A_IWL<9392> A_IWL<9391> A_IWL<9390> A_IWL<9389> A_IWL<9388> A_IWL<9387> A_IWL<9386> A_IWL<9385> A_IWL<9384> A_IWL<9383> A_IWL<9382> A_IWL<9381> A_IWL<9380> A_IWL<9379> A_IWL<9378> A_IWL<9377> A_IWL<9376> A_IWL<9375> A_IWL<9374> A_IWL<9373> A_IWL<9372> A_IWL<9371> A_IWL<9370> A_IWL<9369> A_IWL<9368> A_IWL<9367> A_IWL<9366> A_IWL<9365> A_IWL<9364> A_IWL<9363> A_IWL<9362> A_IWL<9361> A_IWL<9360> A_IWL<9359> A_IWL<9358> A_IWL<9357> A_IWL<9356> A_IWL<9355> A_IWL<9354> A_IWL<9353> A_IWL<9352> A_IWL<9351> A_IWL<9350> A_IWL<9349> A_IWL<9348> A_IWL<9347> A_IWL<9346> A_IWL<9345> A_IWL<9344> A_IWL<9343> A_IWL<9342> A_IWL<9341> A_IWL<9340> A_IWL<9339> A_IWL<9338> A_IWL<9337> A_IWL<9336> A_IWL<9335> A_IWL<9334> A_IWL<9333> A_IWL<9332> A_IWL<9331> A_IWL<9330> A_IWL<9329> A_IWL<9328> A_IWL<9327> A_IWL<9326> A_IWL<9325> A_IWL<9324> A_IWL<9323> A_IWL<9322> A_IWL<9321> A_IWL<9320> A_IWL<9319> A_IWL<9318> A_IWL<9317> A_IWL<9316> A_IWL<9315> A_IWL<9314> A_IWL<9313> A_IWL<9312> A_IWL<9311> A_IWL<9310> A_IWL<9309> A_IWL<9308> A_IWL<9307> A_IWL<9306> A_IWL<9305> A_IWL<9304> A_IWL<9303> A_IWL<9302> A_IWL<9301> A_IWL<9300> A_IWL<9299> A_IWL<9298> A_IWL<9297> A_IWL<9296> A_IWL<9295> A_IWL<9294> A_IWL<9293> A_IWL<9292> A_IWL<9291> A_IWL<9290> A_IWL<9289> A_IWL<9288> A_IWL<9287> A_IWL<9286> A_IWL<9285> A_IWL<9284> A_IWL<9283> A_IWL<9282> A_IWL<9281> A_IWL<9280> A_IWL<9279> A_IWL<9278> A_IWL<9277> A_IWL<9276> A_IWL<9275> A_IWL<9274> A_IWL<9273> A_IWL<9272> A_IWL<9271> A_IWL<9270> A_IWL<9269> A_IWL<9268> A_IWL<9267> A_IWL<9266> A_IWL<9265> A_IWL<9264> A_IWL<9263> A_IWL<9262> A_IWL<9261> A_IWL<9260> A_IWL<9259> A_IWL<9258> A_IWL<9257> A_IWL<9256> A_IWL<9255> A_IWL<9254> A_IWL<9253> A_IWL<9252> A_IWL<9251> A_IWL<9250> A_IWL<9249> A_IWL<9248> A_IWL<9247> A_IWL<9246> A_IWL<9245> A_IWL<9244> A_IWL<9243> A_IWL<9242> A_IWL<9241> A_IWL<9240> A_IWL<9239> A_IWL<9238> A_IWL<9237> A_IWL<9236> A_IWL<9235> A_IWL<9234> A_IWL<9233> A_IWL<9232> A_IWL<9231> A_IWL<9230> A_IWL<9229> A_IWL<9228> A_IWL<9227> A_IWL<9226> A_IWL<9225> A_IWL<9224> A_IWL<9223> A_IWL<9222> A_IWL<9221> A_IWL<9220> A_IWL<9219> A_IWL<9218> A_IWL<9217> A_IWL<9216> A_IWL<9727> A_IWL<9726> A_IWL<9725> A_IWL<9724> A_IWL<9723> A_IWL<9722> A_IWL<9721> A_IWL<9720> A_IWL<9719> A_IWL<9718> A_IWL<9717> A_IWL<9716> A_IWL<9715> A_IWL<9714> A_IWL<9713> A_IWL<9712> A_IWL<9711> A_IWL<9710> A_IWL<9709> A_IWL<9708> A_IWL<9707> A_IWL<9706> A_IWL<9705> A_IWL<9704> A_IWL<9703> A_IWL<9702> A_IWL<9701> A_IWL<9700> A_IWL<9699> A_IWL<9698> A_IWL<9697> A_IWL<9696> A_IWL<9695> A_IWL<9694> A_IWL<9693> A_IWL<9692> A_IWL<9691> A_IWL<9690> A_IWL<9689> A_IWL<9688> A_IWL<9687> A_IWL<9686> A_IWL<9685> A_IWL<9684> A_IWL<9683> A_IWL<9682> A_IWL<9681> A_IWL<9680> A_IWL<9679> A_IWL<9678> A_IWL<9677> A_IWL<9676> A_IWL<9675> A_IWL<9674> A_IWL<9673> A_IWL<9672> A_IWL<9671> A_IWL<9670> A_IWL<9669> A_IWL<9668> A_IWL<9667> A_IWL<9666> A_IWL<9665> A_IWL<9664> A_IWL<9663> A_IWL<9662> A_IWL<9661> A_IWL<9660> A_IWL<9659> A_IWL<9658> A_IWL<9657> A_IWL<9656> A_IWL<9655> A_IWL<9654> A_IWL<9653> A_IWL<9652> A_IWL<9651> A_IWL<9650> A_IWL<9649> A_IWL<9648> A_IWL<9647> A_IWL<9646> A_IWL<9645> A_IWL<9644> A_IWL<9643> A_IWL<9642> A_IWL<9641> A_IWL<9640> A_IWL<9639> A_IWL<9638> A_IWL<9637> A_IWL<9636> A_IWL<9635> A_IWL<9634> A_IWL<9633> A_IWL<9632> A_IWL<9631> A_IWL<9630> A_IWL<9629> A_IWL<9628> A_IWL<9627> A_IWL<9626> A_IWL<9625> A_IWL<9624> A_IWL<9623> A_IWL<9622> A_IWL<9621> A_IWL<9620> A_IWL<9619> A_IWL<9618> A_IWL<9617> A_IWL<9616> A_IWL<9615> A_IWL<9614> A_IWL<9613> A_IWL<9612> A_IWL<9611> A_IWL<9610> A_IWL<9609> A_IWL<9608> A_IWL<9607> A_IWL<9606> A_IWL<9605> A_IWL<9604> A_IWL<9603> A_IWL<9602> A_IWL<9601> A_IWL<9600> A_IWL<9599> A_IWL<9598> A_IWL<9597> A_IWL<9596> A_IWL<9595> A_IWL<9594> A_IWL<9593> A_IWL<9592> A_IWL<9591> A_IWL<9590> A_IWL<9589> A_IWL<9588> A_IWL<9587> A_IWL<9586> A_IWL<9585> A_IWL<9584> A_IWL<9583> A_IWL<9582> A_IWL<9581> A_IWL<9580> A_IWL<9579> A_IWL<9578> A_IWL<9577> A_IWL<9576> A_IWL<9575> A_IWL<9574> A_IWL<9573> A_IWL<9572> A_IWL<9571> A_IWL<9570> A_IWL<9569> A_IWL<9568> A_IWL<9567> A_IWL<9566> A_IWL<9565> A_IWL<9564> A_IWL<9563> A_IWL<9562> A_IWL<9561> A_IWL<9560> A_IWL<9559> A_IWL<9558> A_IWL<9557> A_IWL<9556> A_IWL<9555> A_IWL<9554> A_IWL<9553> A_IWL<9552> A_IWL<9551> A_IWL<9550> A_IWL<9549> A_IWL<9548> A_IWL<9547> A_IWL<9546> A_IWL<9545> A_IWL<9544> A_IWL<9543> A_IWL<9542> A_IWL<9541> A_IWL<9540> A_IWL<9539> A_IWL<9538> A_IWL<9537> A_IWL<9536> A_IWL<9535> A_IWL<9534> A_IWL<9533> A_IWL<9532> A_IWL<9531> A_IWL<9530> A_IWL<9529> A_IWL<9528> A_IWL<9527> A_IWL<9526> A_IWL<9525> A_IWL<9524> A_IWL<9523> A_IWL<9522> A_IWL<9521> A_IWL<9520> A_IWL<9519> A_IWL<9518> A_IWL<9517> A_IWL<9516> A_IWL<9515> A_IWL<9514> A_IWL<9513> A_IWL<9512> A_IWL<9511> A_IWL<9510> A_IWL<9509> A_IWL<9508> A_IWL<9507> A_IWL<9506> A_IWL<9505> A_IWL<9504> A_IWL<9503> A_IWL<9502> A_IWL<9501> A_IWL<9500> A_IWL<9499> A_IWL<9498> A_IWL<9497> A_IWL<9496> A_IWL<9495> A_IWL<9494> A_IWL<9493> A_IWL<9492> A_IWL<9491> A_IWL<9490> A_IWL<9489> A_IWL<9488> A_IWL<9487> A_IWL<9486> A_IWL<9485> A_IWL<9484> A_IWL<9483> A_IWL<9482> A_IWL<9481> A_IWL<9480> A_IWL<9479> A_IWL<9478> A_IWL<9477> A_IWL<9476> A_IWL<9475> A_IWL<9474> A_IWL<9473> A_IWL<9472> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<36> A_BLC<73> A_BLC<72> A_BLC_TOP<73> A_BLC_TOP<72> A_BLT<73> A_BLT<72> A_BLT_TOP<73> A_BLT_TOP<72> A_IWL<9215> A_IWL<9214> A_IWL<9213> A_IWL<9212> A_IWL<9211> A_IWL<9210> A_IWL<9209> A_IWL<9208> A_IWL<9207> A_IWL<9206> A_IWL<9205> A_IWL<9204> A_IWL<9203> A_IWL<9202> A_IWL<9201> A_IWL<9200> A_IWL<9199> A_IWL<9198> A_IWL<9197> A_IWL<9196> A_IWL<9195> A_IWL<9194> A_IWL<9193> A_IWL<9192> A_IWL<9191> A_IWL<9190> A_IWL<9189> A_IWL<9188> A_IWL<9187> A_IWL<9186> A_IWL<9185> A_IWL<9184> A_IWL<9183> A_IWL<9182> A_IWL<9181> A_IWL<9180> A_IWL<9179> A_IWL<9178> A_IWL<9177> A_IWL<9176> A_IWL<9175> A_IWL<9174> A_IWL<9173> A_IWL<9172> A_IWL<9171> A_IWL<9170> A_IWL<9169> A_IWL<9168> A_IWL<9167> A_IWL<9166> A_IWL<9165> A_IWL<9164> A_IWL<9163> A_IWL<9162> A_IWL<9161> A_IWL<9160> A_IWL<9159> A_IWL<9158> A_IWL<9157> A_IWL<9156> A_IWL<9155> A_IWL<9154> A_IWL<9153> A_IWL<9152> A_IWL<9151> A_IWL<9150> A_IWL<9149> A_IWL<9148> A_IWL<9147> A_IWL<9146> A_IWL<9145> A_IWL<9144> A_IWL<9143> A_IWL<9142> A_IWL<9141> A_IWL<9140> A_IWL<9139> A_IWL<9138> A_IWL<9137> A_IWL<9136> A_IWL<9135> A_IWL<9134> A_IWL<9133> A_IWL<9132> A_IWL<9131> A_IWL<9130> A_IWL<9129> A_IWL<9128> A_IWL<9127> A_IWL<9126> A_IWL<9125> A_IWL<9124> A_IWL<9123> A_IWL<9122> A_IWL<9121> A_IWL<9120> A_IWL<9119> A_IWL<9118> A_IWL<9117> A_IWL<9116> A_IWL<9115> A_IWL<9114> A_IWL<9113> A_IWL<9112> A_IWL<9111> A_IWL<9110> A_IWL<9109> A_IWL<9108> A_IWL<9107> A_IWL<9106> A_IWL<9105> A_IWL<9104> A_IWL<9103> A_IWL<9102> A_IWL<9101> A_IWL<9100> A_IWL<9099> A_IWL<9098> A_IWL<9097> A_IWL<9096> A_IWL<9095> A_IWL<9094> A_IWL<9093> A_IWL<9092> A_IWL<9091> A_IWL<9090> A_IWL<9089> A_IWL<9088> A_IWL<9087> A_IWL<9086> A_IWL<9085> A_IWL<9084> A_IWL<9083> A_IWL<9082> A_IWL<9081> A_IWL<9080> A_IWL<9079> A_IWL<9078> A_IWL<9077> A_IWL<9076> A_IWL<9075> A_IWL<9074> A_IWL<9073> A_IWL<9072> A_IWL<9071> A_IWL<9070> A_IWL<9069> A_IWL<9068> A_IWL<9067> A_IWL<9066> A_IWL<9065> A_IWL<9064> A_IWL<9063> A_IWL<9062> A_IWL<9061> A_IWL<9060> A_IWL<9059> A_IWL<9058> A_IWL<9057> A_IWL<9056> A_IWL<9055> A_IWL<9054> A_IWL<9053> A_IWL<9052> A_IWL<9051> A_IWL<9050> A_IWL<9049> A_IWL<9048> A_IWL<9047> A_IWL<9046> A_IWL<9045> A_IWL<9044> A_IWL<9043> A_IWL<9042> A_IWL<9041> A_IWL<9040> A_IWL<9039> A_IWL<9038> A_IWL<9037> A_IWL<9036> A_IWL<9035> A_IWL<9034> A_IWL<9033> A_IWL<9032> A_IWL<9031> A_IWL<9030> A_IWL<9029> A_IWL<9028> A_IWL<9027> A_IWL<9026> A_IWL<9025> A_IWL<9024> A_IWL<9023> A_IWL<9022> A_IWL<9021> A_IWL<9020> A_IWL<9019> A_IWL<9018> A_IWL<9017> A_IWL<9016> A_IWL<9015> A_IWL<9014> A_IWL<9013> A_IWL<9012> A_IWL<9011> A_IWL<9010> A_IWL<9009> A_IWL<9008> A_IWL<9007> A_IWL<9006> A_IWL<9005> A_IWL<9004> A_IWL<9003> A_IWL<9002> A_IWL<9001> A_IWL<9000> A_IWL<8999> A_IWL<8998> A_IWL<8997> A_IWL<8996> A_IWL<8995> A_IWL<8994> A_IWL<8993> A_IWL<8992> A_IWL<8991> A_IWL<8990> A_IWL<8989> A_IWL<8988> A_IWL<8987> A_IWL<8986> A_IWL<8985> A_IWL<8984> A_IWL<8983> A_IWL<8982> A_IWL<8981> A_IWL<8980> A_IWL<8979> A_IWL<8978> A_IWL<8977> A_IWL<8976> A_IWL<8975> A_IWL<8974> A_IWL<8973> A_IWL<8972> A_IWL<8971> A_IWL<8970> A_IWL<8969> A_IWL<8968> A_IWL<8967> A_IWL<8966> A_IWL<8965> A_IWL<8964> A_IWL<8963> A_IWL<8962> A_IWL<8961> A_IWL<8960> A_IWL<9471> A_IWL<9470> A_IWL<9469> A_IWL<9468> A_IWL<9467> A_IWL<9466> A_IWL<9465> A_IWL<9464> A_IWL<9463> A_IWL<9462> A_IWL<9461> A_IWL<9460> A_IWL<9459> A_IWL<9458> A_IWL<9457> A_IWL<9456> A_IWL<9455> A_IWL<9454> A_IWL<9453> A_IWL<9452> A_IWL<9451> A_IWL<9450> A_IWL<9449> A_IWL<9448> A_IWL<9447> A_IWL<9446> A_IWL<9445> A_IWL<9444> A_IWL<9443> A_IWL<9442> A_IWL<9441> A_IWL<9440> A_IWL<9439> A_IWL<9438> A_IWL<9437> A_IWL<9436> A_IWL<9435> A_IWL<9434> A_IWL<9433> A_IWL<9432> A_IWL<9431> A_IWL<9430> A_IWL<9429> A_IWL<9428> A_IWL<9427> A_IWL<9426> A_IWL<9425> A_IWL<9424> A_IWL<9423> A_IWL<9422> A_IWL<9421> A_IWL<9420> A_IWL<9419> A_IWL<9418> A_IWL<9417> A_IWL<9416> A_IWL<9415> A_IWL<9414> A_IWL<9413> A_IWL<9412> A_IWL<9411> A_IWL<9410> A_IWL<9409> A_IWL<9408> A_IWL<9407> A_IWL<9406> A_IWL<9405> A_IWL<9404> A_IWL<9403> A_IWL<9402> A_IWL<9401> A_IWL<9400> A_IWL<9399> A_IWL<9398> A_IWL<9397> A_IWL<9396> A_IWL<9395> A_IWL<9394> A_IWL<9393> A_IWL<9392> A_IWL<9391> A_IWL<9390> A_IWL<9389> A_IWL<9388> A_IWL<9387> A_IWL<9386> A_IWL<9385> A_IWL<9384> A_IWL<9383> A_IWL<9382> A_IWL<9381> A_IWL<9380> A_IWL<9379> A_IWL<9378> A_IWL<9377> A_IWL<9376> A_IWL<9375> A_IWL<9374> A_IWL<9373> A_IWL<9372> A_IWL<9371> A_IWL<9370> A_IWL<9369> A_IWL<9368> A_IWL<9367> A_IWL<9366> A_IWL<9365> A_IWL<9364> A_IWL<9363> A_IWL<9362> A_IWL<9361> A_IWL<9360> A_IWL<9359> A_IWL<9358> A_IWL<9357> A_IWL<9356> A_IWL<9355> A_IWL<9354> A_IWL<9353> A_IWL<9352> A_IWL<9351> A_IWL<9350> A_IWL<9349> A_IWL<9348> A_IWL<9347> A_IWL<9346> A_IWL<9345> A_IWL<9344> A_IWL<9343> A_IWL<9342> A_IWL<9341> A_IWL<9340> A_IWL<9339> A_IWL<9338> A_IWL<9337> A_IWL<9336> A_IWL<9335> A_IWL<9334> A_IWL<9333> A_IWL<9332> A_IWL<9331> A_IWL<9330> A_IWL<9329> A_IWL<9328> A_IWL<9327> A_IWL<9326> A_IWL<9325> A_IWL<9324> A_IWL<9323> A_IWL<9322> A_IWL<9321> A_IWL<9320> A_IWL<9319> A_IWL<9318> A_IWL<9317> A_IWL<9316> A_IWL<9315> A_IWL<9314> A_IWL<9313> A_IWL<9312> A_IWL<9311> A_IWL<9310> A_IWL<9309> A_IWL<9308> A_IWL<9307> A_IWL<9306> A_IWL<9305> A_IWL<9304> A_IWL<9303> A_IWL<9302> A_IWL<9301> A_IWL<9300> A_IWL<9299> A_IWL<9298> A_IWL<9297> A_IWL<9296> A_IWL<9295> A_IWL<9294> A_IWL<9293> A_IWL<9292> A_IWL<9291> A_IWL<9290> A_IWL<9289> A_IWL<9288> A_IWL<9287> A_IWL<9286> A_IWL<9285> A_IWL<9284> A_IWL<9283> A_IWL<9282> A_IWL<9281> A_IWL<9280> A_IWL<9279> A_IWL<9278> A_IWL<9277> A_IWL<9276> A_IWL<9275> A_IWL<9274> A_IWL<9273> A_IWL<9272> A_IWL<9271> A_IWL<9270> A_IWL<9269> A_IWL<9268> A_IWL<9267> A_IWL<9266> A_IWL<9265> A_IWL<9264> A_IWL<9263> A_IWL<9262> A_IWL<9261> A_IWL<9260> A_IWL<9259> A_IWL<9258> A_IWL<9257> A_IWL<9256> A_IWL<9255> A_IWL<9254> A_IWL<9253> A_IWL<9252> A_IWL<9251> A_IWL<9250> A_IWL<9249> A_IWL<9248> A_IWL<9247> A_IWL<9246> A_IWL<9245> A_IWL<9244> A_IWL<9243> A_IWL<9242> A_IWL<9241> A_IWL<9240> A_IWL<9239> A_IWL<9238> A_IWL<9237> A_IWL<9236> A_IWL<9235> A_IWL<9234> A_IWL<9233> A_IWL<9232> A_IWL<9231> A_IWL<9230> A_IWL<9229> A_IWL<9228> A_IWL<9227> A_IWL<9226> A_IWL<9225> A_IWL<9224> A_IWL<9223> A_IWL<9222> A_IWL<9221> A_IWL<9220> A_IWL<9219> A_IWL<9218> A_IWL<9217> A_IWL<9216> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<35> A_BLC<71> A_BLC<70> A_BLC_TOP<71> A_BLC_TOP<70> A_BLT<71> A_BLT<70> A_BLT_TOP<71> A_BLT_TOP<70> A_IWL<8959> A_IWL<8958> A_IWL<8957> A_IWL<8956> A_IWL<8955> A_IWL<8954> A_IWL<8953> A_IWL<8952> A_IWL<8951> A_IWL<8950> A_IWL<8949> A_IWL<8948> A_IWL<8947> A_IWL<8946> A_IWL<8945> A_IWL<8944> A_IWL<8943> A_IWL<8942> A_IWL<8941> A_IWL<8940> A_IWL<8939> A_IWL<8938> A_IWL<8937> A_IWL<8936> A_IWL<8935> A_IWL<8934> A_IWL<8933> A_IWL<8932> A_IWL<8931> A_IWL<8930> A_IWL<8929> A_IWL<8928> A_IWL<8927> A_IWL<8926> A_IWL<8925> A_IWL<8924> A_IWL<8923> A_IWL<8922> A_IWL<8921> A_IWL<8920> A_IWL<8919> A_IWL<8918> A_IWL<8917> A_IWL<8916> A_IWL<8915> A_IWL<8914> A_IWL<8913> A_IWL<8912> A_IWL<8911> A_IWL<8910> A_IWL<8909> A_IWL<8908> A_IWL<8907> A_IWL<8906> A_IWL<8905> A_IWL<8904> A_IWL<8903> A_IWL<8902> A_IWL<8901> A_IWL<8900> A_IWL<8899> A_IWL<8898> A_IWL<8897> A_IWL<8896> A_IWL<8895> A_IWL<8894> A_IWL<8893> A_IWL<8892> A_IWL<8891> A_IWL<8890> A_IWL<8889> A_IWL<8888> A_IWL<8887> A_IWL<8886> A_IWL<8885> A_IWL<8884> A_IWL<8883> A_IWL<8882> A_IWL<8881> A_IWL<8880> A_IWL<8879> A_IWL<8878> A_IWL<8877> A_IWL<8876> A_IWL<8875> A_IWL<8874> A_IWL<8873> A_IWL<8872> A_IWL<8871> A_IWL<8870> A_IWL<8869> A_IWL<8868> A_IWL<8867> A_IWL<8866> A_IWL<8865> A_IWL<8864> A_IWL<8863> A_IWL<8862> A_IWL<8861> A_IWL<8860> A_IWL<8859> A_IWL<8858> A_IWL<8857> A_IWL<8856> A_IWL<8855> A_IWL<8854> A_IWL<8853> A_IWL<8852> A_IWL<8851> A_IWL<8850> A_IWL<8849> A_IWL<8848> A_IWL<8847> A_IWL<8846> A_IWL<8845> A_IWL<8844> A_IWL<8843> A_IWL<8842> A_IWL<8841> A_IWL<8840> A_IWL<8839> A_IWL<8838> A_IWL<8837> A_IWL<8836> A_IWL<8835> A_IWL<8834> A_IWL<8833> A_IWL<8832> A_IWL<8831> A_IWL<8830> A_IWL<8829> A_IWL<8828> A_IWL<8827> A_IWL<8826> A_IWL<8825> A_IWL<8824> A_IWL<8823> A_IWL<8822> A_IWL<8821> A_IWL<8820> A_IWL<8819> A_IWL<8818> A_IWL<8817> A_IWL<8816> A_IWL<8815> A_IWL<8814> A_IWL<8813> A_IWL<8812> A_IWL<8811> A_IWL<8810> A_IWL<8809> A_IWL<8808> A_IWL<8807> A_IWL<8806> A_IWL<8805> A_IWL<8804> A_IWL<8803> A_IWL<8802> A_IWL<8801> A_IWL<8800> A_IWL<8799> A_IWL<8798> A_IWL<8797> A_IWL<8796> A_IWL<8795> A_IWL<8794> A_IWL<8793> A_IWL<8792> A_IWL<8791> A_IWL<8790> A_IWL<8789> A_IWL<8788> A_IWL<8787> A_IWL<8786> A_IWL<8785> A_IWL<8784> A_IWL<8783> A_IWL<8782> A_IWL<8781> A_IWL<8780> A_IWL<8779> A_IWL<8778> A_IWL<8777> A_IWL<8776> A_IWL<8775> A_IWL<8774> A_IWL<8773> A_IWL<8772> A_IWL<8771> A_IWL<8770> A_IWL<8769> A_IWL<8768> A_IWL<8767> A_IWL<8766> A_IWL<8765> A_IWL<8764> A_IWL<8763> A_IWL<8762> A_IWL<8761> A_IWL<8760> A_IWL<8759> A_IWL<8758> A_IWL<8757> A_IWL<8756> A_IWL<8755> A_IWL<8754> A_IWL<8753> A_IWL<8752> A_IWL<8751> A_IWL<8750> A_IWL<8749> A_IWL<8748> A_IWL<8747> A_IWL<8746> A_IWL<8745> A_IWL<8744> A_IWL<8743> A_IWL<8742> A_IWL<8741> A_IWL<8740> A_IWL<8739> A_IWL<8738> A_IWL<8737> A_IWL<8736> A_IWL<8735> A_IWL<8734> A_IWL<8733> A_IWL<8732> A_IWL<8731> A_IWL<8730> A_IWL<8729> A_IWL<8728> A_IWL<8727> A_IWL<8726> A_IWL<8725> A_IWL<8724> A_IWL<8723> A_IWL<8722> A_IWL<8721> A_IWL<8720> A_IWL<8719> A_IWL<8718> A_IWL<8717> A_IWL<8716> A_IWL<8715> A_IWL<8714> A_IWL<8713> A_IWL<8712> A_IWL<8711> A_IWL<8710> A_IWL<8709> A_IWL<8708> A_IWL<8707> A_IWL<8706> A_IWL<8705> A_IWL<8704> A_IWL<9215> A_IWL<9214> A_IWL<9213> A_IWL<9212> A_IWL<9211> A_IWL<9210> A_IWL<9209> A_IWL<9208> A_IWL<9207> A_IWL<9206> A_IWL<9205> A_IWL<9204> A_IWL<9203> A_IWL<9202> A_IWL<9201> A_IWL<9200> A_IWL<9199> A_IWL<9198> A_IWL<9197> A_IWL<9196> A_IWL<9195> A_IWL<9194> A_IWL<9193> A_IWL<9192> A_IWL<9191> A_IWL<9190> A_IWL<9189> A_IWL<9188> A_IWL<9187> A_IWL<9186> A_IWL<9185> A_IWL<9184> A_IWL<9183> A_IWL<9182> A_IWL<9181> A_IWL<9180> A_IWL<9179> A_IWL<9178> A_IWL<9177> A_IWL<9176> A_IWL<9175> A_IWL<9174> A_IWL<9173> A_IWL<9172> A_IWL<9171> A_IWL<9170> A_IWL<9169> A_IWL<9168> A_IWL<9167> A_IWL<9166> A_IWL<9165> A_IWL<9164> A_IWL<9163> A_IWL<9162> A_IWL<9161> A_IWL<9160> A_IWL<9159> A_IWL<9158> A_IWL<9157> A_IWL<9156> A_IWL<9155> A_IWL<9154> A_IWL<9153> A_IWL<9152> A_IWL<9151> A_IWL<9150> A_IWL<9149> A_IWL<9148> A_IWL<9147> A_IWL<9146> A_IWL<9145> A_IWL<9144> A_IWL<9143> A_IWL<9142> A_IWL<9141> A_IWL<9140> A_IWL<9139> A_IWL<9138> A_IWL<9137> A_IWL<9136> A_IWL<9135> A_IWL<9134> A_IWL<9133> A_IWL<9132> A_IWL<9131> A_IWL<9130> A_IWL<9129> A_IWL<9128> A_IWL<9127> A_IWL<9126> A_IWL<9125> A_IWL<9124> A_IWL<9123> A_IWL<9122> A_IWL<9121> A_IWL<9120> A_IWL<9119> A_IWL<9118> A_IWL<9117> A_IWL<9116> A_IWL<9115> A_IWL<9114> A_IWL<9113> A_IWL<9112> A_IWL<9111> A_IWL<9110> A_IWL<9109> A_IWL<9108> A_IWL<9107> A_IWL<9106> A_IWL<9105> A_IWL<9104> A_IWL<9103> A_IWL<9102> A_IWL<9101> A_IWL<9100> A_IWL<9099> A_IWL<9098> A_IWL<9097> A_IWL<9096> A_IWL<9095> A_IWL<9094> A_IWL<9093> A_IWL<9092> A_IWL<9091> A_IWL<9090> A_IWL<9089> A_IWL<9088> A_IWL<9087> A_IWL<9086> A_IWL<9085> A_IWL<9084> A_IWL<9083> A_IWL<9082> A_IWL<9081> A_IWL<9080> A_IWL<9079> A_IWL<9078> A_IWL<9077> A_IWL<9076> A_IWL<9075> A_IWL<9074> A_IWL<9073> A_IWL<9072> A_IWL<9071> A_IWL<9070> A_IWL<9069> A_IWL<9068> A_IWL<9067> A_IWL<9066> A_IWL<9065> A_IWL<9064> A_IWL<9063> A_IWL<9062> A_IWL<9061> A_IWL<9060> A_IWL<9059> A_IWL<9058> A_IWL<9057> A_IWL<9056> A_IWL<9055> A_IWL<9054> A_IWL<9053> A_IWL<9052> A_IWL<9051> A_IWL<9050> A_IWL<9049> A_IWL<9048> A_IWL<9047> A_IWL<9046> A_IWL<9045> A_IWL<9044> A_IWL<9043> A_IWL<9042> A_IWL<9041> A_IWL<9040> A_IWL<9039> A_IWL<9038> A_IWL<9037> A_IWL<9036> A_IWL<9035> A_IWL<9034> A_IWL<9033> A_IWL<9032> A_IWL<9031> A_IWL<9030> A_IWL<9029> A_IWL<9028> A_IWL<9027> A_IWL<9026> A_IWL<9025> A_IWL<9024> A_IWL<9023> A_IWL<9022> A_IWL<9021> A_IWL<9020> A_IWL<9019> A_IWL<9018> A_IWL<9017> A_IWL<9016> A_IWL<9015> A_IWL<9014> A_IWL<9013> A_IWL<9012> A_IWL<9011> A_IWL<9010> A_IWL<9009> A_IWL<9008> A_IWL<9007> A_IWL<9006> A_IWL<9005> A_IWL<9004> A_IWL<9003> A_IWL<9002> A_IWL<9001> A_IWL<9000> A_IWL<8999> A_IWL<8998> A_IWL<8997> A_IWL<8996> A_IWL<8995> A_IWL<8994> A_IWL<8993> A_IWL<8992> A_IWL<8991> A_IWL<8990> A_IWL<8989> A_IWL<8988> A_IWL<8987> A_IWL<8986> A_IWL<8985> A_IWL<8984> A_IWL<8983> A_IWL<8982> A_IWL<8981> A_IWL<8980> A_IWL<8979> A_IWL<8978> A_IWL<8977> A_IWL<8976> A_IWL<8975> A_IWL<8974> A_IWL<8973> A_IWL<8972> A_IWL<8971> A_IWL<8970> A_IWL<8969> A_IWL<8968> A_IWL<8967> A_IWL<8966> A_IWL<8965> A_IWL<8964> A_IWL<8963> A_IWL<8962> A_IWL<8961> A_IWL<8960> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<34> A_BLC<69> A_BLC<68> A_BLC_TOP<69> A_BLC_TOP<68> A_BLT<69> A_BLT<68> A_BLT_TOP<69> A_BLT_TOP<68> A_IWL<8703> A_IWL<8702> A_IWL<8701> A_IWL<8700> A_IWL<8699> A_IWL<8698> A_IWL<8697> A_IWL<8696> A_IWL<8695> A_IWL<8694> A_IWL<8693> A_IWL<8692> A_IWL<8691> A_IWL<8690> A_IWL<8689> A_IWL<8688> A_IWL<8687> A_IWL<8686> A_IWL<8685> A_IWL<8684> A_IWL<8683> A_IWL<8682> A_IWL<8681> A_IWL<8680> A_IWL<8679> A_IWL<8678> A_IWL<8677> A_IWL<8676> A_IWL<8675> A_IWL<8674> A_IWL<8673> A_IWL<8672> A_IWL<8671> A_IWL<8670> A_IWL<8669> A_IWL<8668> A_IWL<8667> A_IWL<8666> A_IWL<8665> A_IWL<8664> A_IWL<8663> A_IWL<8662> A_IWL<8661> A_IWL<8660> A_IWL<8659> A_IWL<8658> A_IWL<8657> A_IWL<8656> A_IWL<8655> A_IWL<8654> A_IWL<8653> A_IWL<8652> A_IWL<8651> A_IWL<8650> A_IWL<8649> A_IWL<8648> A_IWL<8647> A_IWL<8646> A_IWL<8645> A_IWL<8644> A_IWL<8643> A_IWL<8642> A_IWL<8641> A_IWL<8640> A_IWL<8639> A_IWL<8638> A_IWL<8637> A_IWL<8636> A_IWL<8635> A_IWL<8634> A_IWL<8633> A_IWL<8632> A_IWL<8631> A_IWL<8630> A_IWL<8629> A_IWL<8628> A_IWL<8627> A_IWL<8626> A_IWL<8625> A_IWL<8624> A_IWL<8623> A_IWL<8622> A_IWL<8621> A_IWL<8620> A_IWL<8619> A_IWL<8618> A_IWL<8617> A_IWL<8616> A_IWL<8615> A_IWL<8614> A_IWL<8613> A_IWL<8612> A_IWL<8611> A_IWL<8610> A_IWL<8609> A_IWL<8608> A_IWL<8607> A_IWL<8606> A_IWL<8605> A_IWL<8604> A_IWL<8603> A_IWL<8602> A_IWL<8601> A_IWL<8600> A_IWL<8599> A_IWL<8598> A_IWL<8597> A_IWL<8596> A_IWL<8595> A_IWL<8594> A_IWL<8593> A_IWL<8592> A_IWL<8591> A_IWL<8590> A_IWL<8589> A_IWL<8588> A_IWL<8587> A_IWL<8586> A_IWL<8585> A_IWL<8584> A_IWL<8583> A_IWL<8582> A_IWL<8581> A_IWL<8580> A_IWL<8579> A_IWL<8578> A_IWL<8577> A_IWL<8576> A_IWL<8575> A_IWL<8574> A_IWL<8573> A_IWL<8572> A_IWL<8571> A_IWL<8570> A_IWL<8569> A_IWL<8568> A_IWL<8567> A_IWL<8566> A_IWL<8565> A_IWL<8564> A_IWL<8563> A_IWL<8562> A_IWL<8561> A_IWL<8560> A_IWL<8559> A_IWL<8558> A_IWL<8557> A_IWL<8556> A_IWL<8555> A_IWL<8554> A_IWL<8553> A_IWL<8552> A_IWL<8551> A_IWL<8550> A_IWL<8549> A_IWL<8548> A_IWL<8547> A_IWL<8546> A_IWL<8545> A_IWL<8544> A_IWL<8543> A_IWL<8542> A_IWL<8541> A_IWL<8540> A_IWL<8539> A_IWL<8538> A_IWL<8537> A_IWL<8536> A_IWL<8535> A_IWL<8534> A_IWL<8533> A_IWL<8532> A_IWL<8531> A_IWL<8530> A_IWL<8529> A_IWL<8528> A_IWL<8527> A_IWL<8526> A_IWL<8525> A_IWL<8524> A_IWL<8523> A_IWL<8522> A_IWL<8521> A_IWL<8520> A_IWL<8519> A_IWL<8518> A_IWL<8517> A_IWL<8516> A_IWL<8515> A_IWL<8514> A_IWL<8513> A_IWL<8512> A_IWL<8511> A_IWL<8510> A_IWL<8509> A_IWL<8508> A_IWL<8507> A_IWL<8506> A_IWL<8505> A_IWL<8504> A_IWL<8503> A_IWL<8502> A_IWL<8501> A_IWL<8500> A_IWL<8499> A_IWL<8498> A_IWL<8497> A_IWL<8496> A_IWL<8495> A_IWL<8494> A_IWL<8493> A_IWL<8492> A_IWL<8491> A_IWL<8490> A_IWL<8489> A_IWL<8488> A_IWL<8487> A_IWL<8486> A_IWL<8485> A_IWL<8484> A_IWL<8483> A_IWL<8482> A_IWL<8481> A_IWL<8480> A_IWL<8479> A_IWL<8478> A_IWL<8477> A_IWL<8476> A_IWL<8475> A_IWL<8474> A_IWL<8473> A_IWL<8472> A_IWL<8471> A_IWL<8470> A_IWL<8469> A_IWL<8468> A_IWL<8467> A_IWL<8466> A_IWL<8465> A_IWL<8464> A_IWL<8463> A_IWL<8462> A_IWL<8461> A_IWL<8460> A_IWL<8459> A_IWL<8458> A_IWL<8457> A_IWL<8456> A_IWL<8455> A_IWL<8454> A_IWL<8453> A_IWL<8452> A_IWL<8451> A_IWL<8450> A_IWL<8449> A_IWL<8448> A_IWL<8959> A_IWL<8958> A_IWL<8957> A_IWL<8956> A_IWL<8955> A_IWL<8954> A_IWL<8953> A_IWL<8952> A_IWL<8951> A_IWL<8950> A_IWL<8949> A_IWL<8948> A_IWL<8947> A_IWL<8946> A_IWL<8945> A_IWL<8944> A_IWL<8943> A_IWL<8942> A_IWL<8941> A_IWL<8940> A_IWL<8939> A_IWL<8938> A_IWL<8937> A_IWL<8936> A_IWL<8935> A_IWL<8934> A_IWL<8933> A_IWL<8932> A_IWL<8931> A_IWL<8930> A_IWL<8929> A_IWL<8928> A_IWL<8927> A_IWL<8926> A_IWL<8925> A_IWL<8924> A_IWL<8923> A_IWL<8922> A_IWL<8921> A_IWL<8920> A_IWL<8919> A_IWL<8918> A_IWL<8917> A_IWL<8916> A_IWL<8915> A_IWL<8914> A_IWL<8913> A_IWL<8912> A_IWL<8911> A_IWL<8910> A_IWL<8909> A_IWL<8908> A_IWL<8907> A_IWL<8906> A_IWL<8905> A_IWL<8904> A_IWL<8903> A_IWL<8902> A_IWL<8901> A_IWL<8900> A_IWL<8899> A_IWL<8898> A_IWL<8897> A_IWL<8896> A_IWL<8895> A_IWL<8894> A_IWL<8893> A_IWL<8892> A_IWL<8891> A_IWL<8890> A_IWL<8889> A_IWL<8888> A_IWL<8887> A_IWL<8886> A_IWL<8885> A_IWL<8884> A_IWL<8883> A_IWL<8882> A_IWL<8881> A_IWL<8880> A_IWL<8879> A_IWL<8878> A_IWL<8877> A_IWL<8876> A_IWL<8875> A_IWL<8874> A_IWL<8873> A_IWL<8872> A_IWL<8871> A_IWL<8870> A_IWL<8869> A_IWL<8868> A_IWL<8867> A_IWL<8866> A_IWL<8865> A_IWL<8864> A_IWL<8863> A_IWL<8862> A_IWL<8861> A_IWL<8860> A_IWL<8859> A_IWL<8858> A_IWL<8857> A_IWL<8856> A_IWL<8855> A_IWL<8854> A_IWL<8853> A_IWL<8852> A_IWL<8851> A_IWL<8850> A_IWL<8849> A_IWL<8848> A_IWL<8847> A_IWL<8846> A_IWL<8845> A_IWL<8844> A_IWL<8843> A_IWL<8842> A_IWL<8841> A_IWL<8840> A_IWL<8839> A_IWL<8838> A_IWL<8837> A_IWL<8836> A_IWL<8835> A_IWL<8834> A_IWL<8833> A_IWL<8832> A_IWL<8831> A_IWL<8830> A_IWL<8829> A_IWL<8828> A_IWL<8827> A_IWL<8826> A_IWL<8825> A_IWL<8824> A_IWL<8823> A_IWL<8822> A_IWL<8821> A_IWL<8820> A_IWL<8819> A_IWL<8818> A_IWL<8817> A_IWL<8816> A_IWL<8815> A_IWL<8814> A_IWL<8813> A_IWL<8812> A_IWL<8811> A_IWL<8810> A_IWL<8809> A_IWL<8808> A_IWL<8807> A_IWL<8806> A_IWL<8805> A_IWL<8804> A_IWL<8803> A_IWL<8802> A_IWL<8801> A_IWL<8800> A_IWL<8799> A_IWL<8798> A_IWL<8797> A_IWL<8796> A_IWL<8795> A_IWL<8794> A_IWL<8793> A_IWL<8792> A_IWL<8791> A_IWL<8790> A_IWL<8789> A_IWL<8788> A_IWL<8787> A_IWL<8786> A_IWL<8785> A_IWL<8784> A_IWL<8783> A_IWL<8782> A_IWL<8781> A_IWL<8780> A_IWL<8779> A_IWL<8778> A_IWL<8777> A_IWL<8776> A_IWL<8775> A_IWL<8774> A_IWL<8773> A_IWL<8772> A_IWL<8771> A_IWL<8770> A_IWL<8769> A_IWL<8768> A_IWL<8767> A_IWL<8766> A_IWL<8765> A_IWL<8764> A_IWL<8763> A_IWL<8762> A_IWL<8761> A_IWL<8760> A_IWL<8759> A_IWL<8758> A_IWL<8757> A_IWL<8756> A_IWL<8755> A_IWL<8754> A_IWL<8753> A_IWL<8752> A_IWL<8751> A_IWL<8750> A_IWL<8749> A_IWL<8748> A_IWL<8747> A_IWL<8746> A_IWL<8745> A_IWL<8744> A_IWL<8743> A_IWL<8742> A_IWL<8741> A_IWL<8740> A_IWL<8739> A_IWL<8738> A_IWL<8737> A_IWL<8736> A_IWL<8735> A_IWL<8734> A_IWL<8733> A_IWL<8732> A_IWL<8731> A_IWL<8730> A_IWL<8729> A_IWL<8728> A_IWL<8727> A_IWL<8726> A_IWL<8725> A_IWL<8724> A_IWL<8723> A_IWL<8722> A_IWL<8721> A_IWL<8720> A_IWL<8719> A_IWL<8718> A_IWL<8717> A_IWL<8716> A_IWL<8715> A_IWL<8714> A_IWL<8713> A_IWL<8712> A_IWL<8711> A_IWL<8710> A_IWL<8709> A_IWL<8708> A_IWL<8707> A_IWL<8706> A_IWL<8705> A_IWL<8704> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<33> A_BLC<67> A_BLC<66> A_BLC_TOP<67> A_BLC_TOP<66> A_BLT<67> A_BLT<66> A_BLT_TOP<67> A_BLT_TOP<66> A_IWL<8447> A_IWL<8446> A_IWL<8445> A_IWL<8444> A_IWL<8443> A_IWL<8442> A_IWL<8441> A_IWL<8440> A_IWL<8439> A_IWL<8438> A_IWL<8437> A_IWL<8436> A_IWL<8435> A_IWL<8434> A_IWL<8433> A_IWL<8432> A_IWL<8431> A_IWL<8430> A_IWL<8429> A_IWL<8428> A_IWL<8427> A_IWL<8426> A_IWL<8425> A_IWL<8424> A_IWL<8423> A_IWL<8422> A_IWL<8421> A_IWL<8420> A_IWL<8419> A_IWL<8418> A_IWL<8417> A_IWL<8416> A_IWL<8415> A_IWL<8414> A_IWL<8413> A_IWL<8412> A_IWL<8411> A_IWL<8410> A_IWL<8409> A_IWL<8408> A_IWL<8407> A_IWL<8406> A_IWL<8405> A_IWL<8404> A_IWL<8403> A_IWL<8402> A_IWL<8401> A_IWL<8400> A_IWL<8399> A_IWL<8398> A_IWL<8397> A_IWL<8396> A_IWL<8395> A_IWL<8394> A_IWL<8393> A_IWL<8392> A_IWL<8391> A_IWL<8390> A_IWL<8389> A_IWL<8388> A_IWL<8387> A_IWL<8386> A_IWL<8385> A_IWL<8384> A_IWL<8383> A_IWL<8382> A_IWL<8381> A_IWL<8380> A_IWL<8379> A_IWL<8378> A_IWL<8377> A_IWL<8376> A_IWL<8375> A_IWL<8374> A_IWL<8373> A_IWL<8372> A_IWL<8371> A_IWL<8370> A_IWL<8369> A_IWL<8368> A_IWL<8367> A_IWL<8366> A_IWL<8365> A_IWL<8364> A_IWL<8363> A_IWL<8362> A_IWL<8361> A_IWL<8360> A_IWL<8359> A_IWL<8358> A_IWL<8357> A_IWL<8356> A_IWL<8355> A_IWL<8354> A_IWL<8353> A_IWL<8352> A_IWL<8351> A_IWL<8350> A_IWL<8349> A_IWL<8348> A_IWL<8347> A_IWL<8346> A_IWL<8345> A_IWL<8344> A_IWL<8343> A_IWL<8342> A_IWL<8341> A_IWL<8340> A_IWL<8339> A_IWL<8338> A_IWL<8337> A_IWL<8336> A_IWL<8335> A_IWL<8334> A_IWL<8333> A_IWL<8332> A_IWL<8331> A_IWL<8330> A_IWL<8329> A_IWL<8328> A_IWL<8327> A_IWL<8326> A_IWL<8325> A_IWL<8324> A_IWL<8323> A_IWL<8322> A_IWL<8321> A_IWL<8320> A_IWL<8319> A_IWL<8318> A_IWL<8317> A_IWL<8316> A_IWL<8315> A_IWL<8314> A_IWL<8313> A_IWL<8312> A_IWL<8311> A_IWL<8310> A_IWL<8309> A_IWL<8308> A_IWL<8307> A_IWL<8306> A_IWL<8305> A_IWL<8304> A_IWL<8303> A_IWL<8302> A_IWL<8301> A_IWL<8300> A_IWL<8299> A_IWL<8298> A_IWL<8297> A_IWL<8296> A_IWL<8295> A_IWL<8294> A_IWL<8293> A_IWL<8292> A_IWL<8291> A_IWL<8290> A_IWL<8289> A_IWL<8288> A_IWL<8287> A_IWL<8286> A_IWL<8285> A_IWL<8284> A_IWL<8283> A_IWL<8282> A_IWL<8281> A_IWL<8280> A_IWL<8279> A_IWL<8278> A_IWL<8277> A_IWL<8276> A_IWL<8275> A_IWL<8274> A_IWL<8273> A_IWL<8272> A_IWL<8271> A_IWL<8270> A_IWL<8269> A_IWL<8268> A_IWL<8267> A_IWL<8266> A_IWL<8265> A_IWL<8264> A_IWL<8263> A_IWL<8262> A_IWL<8261> A_IWL<8260> A_IWL<8259> A_IWL<8258> A_IWL<8257> A_IWL<8256> A_IWL<8255> A_IWL<8254> A_IWL<8253> A_IWL<8252> A_IWL<8251> A_IWL<8250> A_IWL<8249> A_IWL<8248> A_IWL<8247> A_IWL<8246> A_IWL<8245> A_IWL<8244> A_IWL<8243> A_IWL<8242> A_IWL<8241> A_IWL<8240> A_IWL<8239> A_IWL<8238> A_IWL<8237> A_IWL<8236> A_IWL<8235> A_IWL<8234> A_IWL<8233> A_IWL<8232> A_IWL<8231> A_IWL<8230> A_IWL<8229> A_IWL<8228> A_IWL<8227> A_IWL<8226> A_IWL<8225> A_IWL<8224> A_IWL<8223> A_IWL<8222> A_IWL<8221> A_IWL<8220> A_IWL<8219> A_IWL<8218> A_IWL<8217> A_IWL<8216> A_IWL<8215> A_IWL<8214> A_IWL<8213> A_IWL<8212> A_IWL<8211> A_IWL<8210> A_IWL<8209> A_IWL<8208> A_IWL<8207> A_IWL<8206> A_IWL<8205> A_IWL<8204> A_IWL<8203> A_IWL<8202> A_IWL<8201> A_IWL<8200> A_IWL<8199> A_IWL<8198> A_IWL<8197> A_IWL<8196> A_IWL<8195> A_IWL<8194> A_IWL<8193> A_IWL<8192> A_IWL<8703> A_IWL<8702> A_IWL<8701> A_IWL<8700> A_IWL<8699> A_IWL<8698> A_IWL<8697> A_IWL<8696> A_IWL<8695> A_IWL<8694> A_IWL<8693> A_IWL<8692> A_IWL<8691> A_IWL<8690> A_IWL<8689> A_IWL<8688> A_IWL<8687> A_IWL<8686> A_IWL<8685> A_IWL<8684> A_IWL<8683> A_IWL<8682> A_IWL<8681> A_IWL<8680> A_IWL<8679> A_IWL<8678> A_IWL<8677> A_IWL<8676> A_IWL<8675> A_IWL<8674> A_IWL<8673> A_IWL<8672> A_IWL<8671> A_IWL<8670> A_IWL<8669> A_IWL<8668> A_IWL<8667> A_IWL<8666> A_IWL<8665> A_IWL<8664> A_IWL<8663> A_IWL<8662> A_IWL<8661> A_IWL<8660> A_IWL<8659> A_IWL<8658> A_IWL<8657> A_IWL<8656> A_IWL<8655> A_IWL<8654> A_IWL<8653> A_IWL<8652> A_IWL<8651> A_IWL<8650> A_IWL<8649> A_IWL<8648> A_IWL<8647> A_IWL<8646> A_IWL<8645> A_IWL<8644> A_IWL<8643> A_IWL<8642> A_IWL<8641> A_IWL<8640> A_IWL<8639> A_IWL<8638> A_IWL<8637> A_IWL<8636> A_IWL<8635> A_IWL<8634> A_IWL<8633> A_IWL<8632> A_IWL<8631> A_IWL<8630> A_IWL<8629> A_IWL<8628> A_IWL<8627> A_IWL<8626> A_IWL<8625> A_IWL<8624> A_IWL<8623> A_IWL<8622> A_IWL<8621> A_IWL<8620> A_IWL<8619> A_IWL<8618> A_IWL<8617> A_IWL<8616> A_IWL<8615> A_IWL<8614> A_IWL<8613> A_IWL<8612> A_IWL<8611> A_IWL<8610> A_IWL<8609> A_IWL<8608> A_IWL<8607> A_IWL<8606> A_IWL<8605> A_IWL<8604> A_IWL<8603> A_IWL<8602> A_IWL<8601> A_IWL<8600> A_IWL<8599> A_IWL<8598> A_IWL<8597> A_IWL<8596> A_IWL<8595> A_IWL<8594> A_IWL<8593> A_IWL<8592> A_IWL<8591> A_IWL<8590> A_IWL<8589> A_IWL<8588> A_IWL<8587> A_IWL<8586> A_IWL<8585> A_IWL<8584> A_IWL<8583> A_IWL<8582> A_IWL<8581> A_IWL<8580> A_IWL<8579> A_IWL<8578> A_IWL<8577> A_IWL<8576> A_IWL<8575> A_IWL<8574> A_IWL<8573> A_IWL<8572> A_IWL<8571> A_IWL<8570> A_IWL<8569> A_IWL<8568> A_IWL<8567> A_IWL<8566> A_IWL<8565> A_IWL<8564> A_IWL<8563> A_IWL<8562> A_IWL<8561> A_IWL<8560> A_IWL<8559> A_IWL<8558> A_IWL<8557> A_IWL<8556> A_IWL<8555> A_IWL<8554> A_IWL<8553> A_IWL<8552> A_IWL<8551> A_IWL<8550> A_IWL<8549> A_IWL<8548> A_IWL<8547> A_IWL<8546> A_IWL<8545> A_IWL<8544> A_IWL<8543> A_IWL<8542> A_IWL<8541> A_IWL<8540> A_IWL<8539> A_IWL<8538> A_IWL<8537> A_IWL<8536> A_IWL<8535> A_IWL<8534> A_IWL<8533> A_IWL<8532> A_IWL<8531> A_IWL<8530> A_IWL<8529> A_IWL<8528> A_IWL<8527> A_IWL<8526> A_IWL<8525> A_IWL<8524> A_IWL<8523> A_IWL<8522> A_IWL<8521> A_IWL<8520> A_IWL<8519> A_IWL<8518> A_IWL<8517> A_IWL<8516> A_IWL<8515> A_IWL<8514> A_IWL<8513> A_IWL<8512> A_IWL<8511> A_IWL<8510> A_IWL<8509> A_IWL<8508> A_IWL<8507> A_IWL<8506> A_IWL<8505> A_IWL<8504> A_IWL<8503> A_IWL<8502> A_IWL<8501> A_IWL<8500> A_IWL<8499> A_IWL<8498> A_IWL<8497> A_IWL<8496> A_IWL<8495> A_IWL<8494> A_IWL<8493> A_IWL<8492> A_IWL<8491> A_IWL<8490> A_IWL<8489> A_IWL<8488> A_IWL<8487> A_IWL<8486> A_IWL<8485> A_IWL<8484> A_IWL<8483> A_IWL<8482> A_IWL<8481> A_IWL<8480> A_IWL<8479> A_IWL<8478> A_IWL<8477> A_IWL<8476> A_IWL<8475> A_IWL<8474> A_IWL<8473> A_IWL<8472> A_IWL<8471> A_IWL<8470> A_IWL<8469> A_IWL<8468> A_IWL<8467> A_IWL<8466> A_IWL<8465> A_IWL<8464> A_IWL<8463> A_IWL<8462> A_IWL<8461> A_IWL<8460> A_IWL<8459> A_IWL<8458> A_IWL<8457> A_IWL<8456> A_IWL<8455> A_IWL<8454> A_IWL<8453> A_IWL<8452> A_IWL<8451> A_IWL<8450> A_IWL<8449> A_IWL<8448> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<32> A_BLC<65> A_BLC<64> A_BLC_TOP<65> A_BLC_TOP<64> A_BLT<65> A_BLT<64> A_BLT_TOP<65> A_BLT_TOP<64> A_IWL<8191> A_IWL<8190> A_IWL<8189> A_IWL<8188> A_IWL<8187> A_IWL<8186> A_IWL<8185> A_IWL<8184> A_IWL<8183> A_IWL<8182> A_IWL<8181> A_IWL<8180> A_IWL<8179> A_IWL<8178> A_IWL<8177> A_IWL<8176> A_IWL<8175> A_IWL<8174> A_IWL<8173> A_IWL<8172> A_IWL<8171> A_IWL<8170> A_IWL<8169> A_IWL<8168> A_IWL<8167> A_IWL<8166> A_IWL<8165> A_IWL<8164> A_IWL<8163> A_IWL<8162> A_IWL<8161> A_IWL<8160> A_IWL<8159> A_IWL<8158> A_IWL<8157> A_IWL<8156> A_IWL<8155> A_IWL<8154> A_IWL<8153> A_IWL<8152> A_IWL<8151> A_IWL<8150> A_IWL<8149> A_IWL<8148> A_IWL<8147> A_IWL<8146> A_IWL<8145> A_IWL<8144> A_IWL<8143> A_IWL<8142> A_IWL<8141> A_IWL<8140> A_IWL<8139> A_IWL<8138> A_IWL<8137> A_IWL<8136> A_IWL<8135> A_IWL<8134> A_IWL<8133> A_IWL<8132> A_IWL<8131> A_IWL<8130> A_IWL<8129> A_IWL<8128> A_IWL<8127> A_IWL<8126> A_IWL<8125> A_IWL<8124> A_IWL<8123> A_IWL<8122> A_IWL<8121> A_IWL<8120> A_IWL<8119> A_IWL<8118> A_IWL<8117> A_IWL<8116> A_IWL<8115> A_IWL<8114> A_IWL<8113> A_IWL<8112> A_IWL<8111> A_IWL<8110> A_IWL<8109> A_IWL<8108> A_IWL<8107> A_IWL<8106> A_IWL<8105> A_IWL<8104> A_IWL<8103> A_IWL<8102> A_IWL<8101> A_IWL<8100> A_IWL<8099> A_IWL<8098> A_IWL<8097> A_IWL<8096> A_IWL<8095> A_IWL<8094> A_IWL<8093> A_IWL<8092> A_IWL<8091> A_IWL<8090> A_IWL<8089> A_IWL<8088> A_IWL<8087> A_IWL<8086> A_IWL<8085> A_IWL<8084> A_IWL<8083> A_IWL<8082> A_IWL<8081> A_IWL<8080> A_IWL<8079> A_IWL<8078> A_IWL<8077> A_IWL<8076> A_IWL<8075> A_IWL<8074> A_IWL<8073> A_IWL<8072> A_IWL<8071> A_IWL<8070> A_IWL<8069> A_IWL<8068> A_IWL<8067> A_IWL<8066> A_IWL<8065> A_IWL<8064> A_IWL<8063> A_IWL<8062> A_IWL<8061> A_IWL<8060> A_IWL<8059> A_IWL<8058> A_IWL<8057> A_IWL<8056> A_IWL<8055> A_IWL<8054> A_IWL<8053> A_IWL<8052> A_IWL<8051> A_IWL<8050> A_IWL<8049> A_IWL<8048> A_IWL<8047> A_IWL<8046> A_IWL<8045> A_IWL<8044> A_IWL<8043> A_IWL<8042> A_IWL<8041> A_IWL<8040> A_IWL<8039> A_IWL<8038> A_IWL<8037> A_IWL<8036> A_IWL<8035> A_IWL<8034> A_IWL<8033> A_IWL<8032> A_IWL<8031> A_IWL<8030> A_IWL<8029> A_IWL<8028> A_IWL<8027> A_IWL<8026> A_IWL<8025> A_IWL<8024> A_IWL<8023> A_IWL<8022> A_IWL<8021> A_IWL<8020> A_IWL<8019> A_IWL<8018> A_IWL<8017> A_IWL<8016> A_IWL<8015> A_IWL<8014> A_IWL<8013> A_IWL<8012> A_IWL<8011> A_IWL<8010> A_IWL<8009> A_IWL<8008> A_IWL<8007> A_IWL<8006> A_IWL<8005> A_IWL<8004> A_IWL<8003> A_IWL<8002> A_IWL<8001> A_IWL<8000> A_IWL<7999> A_IWL<7998> A_IWL<7997> A_IWL<7996> A_IWL<7995> A_IWL<7994> A_IWL<7993> A_IWL<7992> A_IWL<7991> A_IWL<7990> A_IWL<7989> A_IWL<7988> A_IWL<7987> A_IWL<7986> A_IWL<7985> A_IWL<7984> A_IWL<7983> A_IWL<7982> A_IWL<7981> A_IWL<7980> A_IWL<7979> A_IWL<7978> A_IWL<7977> A_IWL<7976> A_IWL<7975> A_IWL<7974> A_IWL<7973> A_IWL<7972> A_IWL<7971> A_IWL<7970> A_IWL<7969> A_IWL<7968> A_IWL<7967> A_IWL<7966> A_IWL<7965> A_IWL<7964> A_IWL<7963> A_IWL<7962> A_IWL<7961> A_IWL<7960> A_IWL<7959> A_IWL<7958> A_IWL<7957> A_IWL<7956> A_IWL<7955> A_IWL<7954> A_IWL<7953> A_IWL<7952> A_IWL<7951> A_IWL<7950> A_IWL<7949> A_IWL<7948> A_IWL<7947> A_IWL<7946> A_IWL<7945> A_IWL<7944> A_IWL<7943> A_IWL<7942> A_IWL<7941> A_IWL<7940> A_IWL<7939> A_IWL<7938> A_IWL<7937> A_IWL<7936> A_IWL<8447> A_IWL<8446> A_IWL<8445> A_IWL<8444> A_IWL<8443> A_IWL<8442> A_IWL<8441> A_IWL<8440> A_IWL<8439> A_IWL<8438> A_IWL<8437> A_IWL<8436> A_IWL<8435> A_IWL<8434> A_IWL<8433> A_IWL<8432> A_IWL<8431> A_IWL<8430> A_IWL<8429> A_IWL<8428> A_IWL<8427> A_IWL<8426> A_IWL<8425> A_IWL<8424> A_IWL<8423> A_IWL<8422> A_IWL<8421> A_IWL<8420> A_IWL<8419> A_IWL<8418> A_IWL<8417> A_IWL<8416> A_IWL<8415> A_IWL<8414> A_IWL<8413> A_IWL<8412> A_IWL<8411> A_IWL<8410> A_IWL<8409> A_IWL<8408> A_IWL<8407> A_IWL<8406> A_IWL<8405> A_IWL<8404> A_IWL<8403> A_IWL<8402> A_IWL<8401> A_IWL<8400> A_IWL<8399> A_IWL<8398> A_IWL<8397> A_IWL<8396> A_IWL<8395> A_IWL<8394> A_IWL<8393> A_IWL<8392> A_IWL<8391> A_IWL<8390> A_IWL<8389> A_IWL<8388> A_IWL<8387> A_IWL<8386> A_IWL<8385> A_IWL<8384> A_IWL<8383> A_IWL<8382> A_IWL<8381> A_IWL<8380> A_IWL<8379> A_IWL<8378> A_IWL<8377> A_IWL<8376> A_IWL<8375> A_IWL<8374> A_IWL<8373> A_IWL<8372> A_IWL<8371> A_IWL<8370> A_IWL<8369> A_IWL<8368> A_IWL<8367> A_IWL<8366> A_IWL<8365> A_IWL<8364> A_IWL<8363> A_IWL<8362> A_IWL<8361> A_IWL<8360> A_IWL<8359> A_IWL<8358> A_IWL<8357> A_IWL<8356> A_IWL<8355> A_IWL<8354> A_IWL<8353> A_IWL<8352> A_IWL<8351> A_IWL<8350> A_IWL<8349> A_IWL<8348> A_IWL<8347> A_IWL<8346> A_IWL<8345> A_IWL<8344> A_IWL<8343> A_IWL<8342> A_IWL<8341> A_IWL<8340> A_IWL<8339> A_IWL<8338> A_IWL<8337> A_IWL<8336> A_IWL<8335> A_IWL<8334> A_IWL<8333> A_IWL<8332> A_IWL<8331> A_IWL<8330> A_IWL<8329> A_IWL<8328> A_IWL<8327> A_IWL<8326> A_IWL<8325> A_IWL<8324> A_IWL<8323> A_IWL<8322> A_IWL<8321> A_IWL<8320> A_IWL<8319> A_IWL<8318> A_IWL<8317> A_IWL<8316> A_IWL<8315> A_IWL<8314> A_IWL<8313> A_IWL<8312> A_IWL<8311> A_IWL<8310> A_IWL<8309> A_IWL<8308> A_IWL<8307> A_IWL<8306> A_IWL<8305> A_IWL<8304> A_IWL<8303> A_IWL<8302> A_IWL<8301> A_IWL<8300> A_IWL<8299> A_IWL<8298> A_IWL<8297> A_IWL<8296> A_IWL<8295> A_IWL<8294> A_IWL<8293> A_IWL<8292> A_IWL<8291> A_IWL<8290> A_IWL<8289> A_IWL<8288> A_IWL<8287> A_IWL<8286> A_IWL<8285> A_IWL<8284> A_IWL<8283> A_IWL<8282> A_IWL<8281> A_IWL<8280> A_IWL<8279> A_IWL<8278> A_IWL<8277> A_IWL<8276> A_IWL<8275> A_IWL<8274> A_IWL<8273> A_IWL<8272> A_IWL<8271> A_IWL<8270> A_IWL<8269> A_IWL<8268> A_IWL<8267> A_IWL<8266> A_IWL<8265> A_IWL<8264> A_IWL<8263> A_IWL<8262> A_IWL<8261> A_IWL<8260> A_IWL<8259> A_IWL<8258> A_IWL<8257> A_IWL<8256> A_IWL<8255> A_IWL<8254> A_IWL<8253> A_IWL<8252> A_IWL<8251> A_IWL<8250> A_IWL<8249> A_IWL<8248> A_IWL<8247> A_IWL<8246> A_IWL<8245> A_IWL<8244> A_IWL<8243> A_IWL<8242> A_IWL<8241> A_IWL<8240> A_IWL<8239> A_IWL<8238> A_IWL<8237> A_IWL<8236> A_IWL<8235> A_IWL<8234> A_IWL<8233> A_IWL<8232> A_IWL<8231> A_IWL<8230> A_IWL<8229> A_IWL<8228> A_IWL<8227> A_IWL<8226> A_IWL<8225> A_IWL<8224> A_IWL<8223> A_IWL<8222> A_IWL<8221> A_IWL<8220> A_IWL<8219> A_IWL<8218> A_IWL<8217> A_IWL<8216> A_IWL<8215> A_IWL<8214> A_IWL<8213> A_IWL<8212> A_IWL<8211> A_IWL<8210> A_IWL<8209> A_IWL<8208> A_IWL<8207> A_IWL<8206> A_IWL<8205> A_IWL<8204> A_IWL<8203> A_IWL<8202> A_IWL<8201> A_IWL<8200> A_IWL<8199> A_IWL<8198> A_IWL<8197> A_IWL<8196> A_IWL<8195> A_IWL<8194> A_IWL<8193> A_IWL<8192> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<31> A_BLC<63> A_BLC<62> A_BLC_TOP<63> A_BLC_TOP<62> A_BLT<63> A_BLT<62> A_BLT_TOP<63> A_BLT_TOP<62> A_IWL<7935> A_IWL<7934> A_IWL<7933> A_IWL<7932> A_IWL<7931> A_IWL<7930> A_IWL<7929> A_IWL<7928> A_IWL<7927> A_IWL<7926> A_IWL<7925> A_IWL<7924> A_IWL<7923> A_IWL<7922> A_IWL<7921> A_IWL<7920> A_IWL<7919> A_IWL<7918> A_IWL<7917> A_IWL<7916> A_IWL<7915> A_IWL<7914> A_IWL<7913> A_IWL<7912> A_IWL<7911> A_IWL<7910> A_IWL<7909> A_IWL<7908> A_IWL<7907> A_IWL<7906> A_IWL<7905> A_IWL<7904> A_IWL<7903> A_IWL<7902> A_IWL<7901> A_IWL<7900> A_IWL<7899> A_IWL<7898> A_IWL<7897> A_IWL<7896> A_IWL<7895> A_IWL<7894> A_IWL<7893> A_IWL<7892> A_IWL<7891> A_IWL<7890> A_IWL<7889> A_IWL<7888> A_IWL<7887> A_IWL<7886> A_IWL<7885> A_IWL<7884> A_IWL<7883> A_IWL<7882> A_IWL<7881> A_IWL<7880> A_IWL<7879> A_IWL<7878> A_IWL<7877> A_IWL<7876> A_IWL<7875> A_IWL<7874> A_IWL<7873> A_IWL<7872> A_IWL<7871> A_IWL<7870> A_IWL<7869> A_IWL<7868> A_IWL<7867> A_IWL<7866> A_IWL<7865> A_IWL<7864> A_IWL<7863> A_IWL<7862> A_IWL<7861> A_IWL<7860> A_IWL<7859> A_IWL<7858> A_IWL<7857> A_IWL<7856> A_IWL<7855> A_IWL<7854> A_IWL<7853> A_IWL<7852> A_IWL<7851> A_IWL<7850> A_IWL<7849> A_IWL<7848> A_IWL<7847> A_IWL<7846> A_IWL<7845> A_IWL<7844> A_IWL<7843> A_IWL<7842> A_IWL<7841> A_IWL<7840> A_IWL<7839> A_IWL<7838> A_IWL<7837> A_IWL<7836> A_IWL<7835> A_IWL<7834> A_IWL<7833> A_IWL<7832> A_IWL<7831> A_IWL<7830> A_IWL<7829> A_IWL<7828> A_IWL<7827> A_IWL<7826> A_IWL<7825> A_IWL<7824> A_IWL<7823> A_IWL<7822> A_IWL<7821> A_IWL<7820> A_IWL<7819> A_IWL<7818> A_IWL<7817> A_IWL<7816> A_IWL<7815> A_IWL<7814> A_IWL<7813> A_IWL<7812> A_IWL<7811> A_IWL<7810> A_IWL<7809> A_IWL<7808> A_IWL<7807> A_IWL<7806> A_IWL<7805> A_IWL<7804> A_IWL<7803> A_IWL<7802> A_IWL<7801> A_IWL<7800> A_IWL<7799> A_IWL<7798> A_IWL<7797> A_IWL<7796> A_IWL<7795> A_IWL<7794> A_IWL<7793> A_IWL<7792> A_IWL<7791> A_IWL<7790> A_IWL<7789> A_IWL<7788> A_IWL<7787> A_IWL<7786> A_IWL<7785> A_IWL<7784> A_IWL<7783> A_IWL<7782> A_IWL<7781> A_IWL<7780> A_IWL<7779> A_IWL<7778> A_IWL<7777> A_IWL<7776> A_IWL<7775> A_IWL<7774> A_IWL<7773> A_IWL<7772> A_IWL<7771> A_IWL<7770> A_IWL<7769> A_IWL<7768> A_IWL<7767> A_IWL<7766> A_IWL<7765> A_IWL<7764> A_IWL<7763> A_IWL<7762> A_IWL<7761> A_IWL<7760> A_IWL<7759> A_IWL<7758> A_IWL<7757> A_IWL<7756> A_IWL<7755> A_IWL<7754> A_IWL<7753> A_IWL<7752> A_IWL<7751> A_IWL<7750> A_IWL<7749> A_IWL<7748> A_IWL<7747> A_IWL<7746> A_IWL<7745> A_IWL<7744> A_IWL<7743> A_IWL<7742> A_IWL<7741> A_IWL<7740> A_IWL<7739> A_IWL<7738> A_IWL<7737> A_IWL<7736> A_IWL<7735> A_IWL<7734> A_IWL<7733> A_IWL<7732> A_IWL<7731> A_IWL<7730> A_IWL<7729> A_IWL<7728> A_IWL<7727> A_IWL<7726> A_IWL<7725> A_IWL<7724> A_IWL<7723> A_IWL<7722> A_IWL<7721> A_IWL<7720> A_IWL<7719> A_IWL<7718> A_IWL<7717> A_IWL<7716> A_IWL<7715> A_IWL<7714> A_IWL<7713> A_IWL<7712> A_IWL<7711> A_IWL<7710> A_IWL<7709> A_IWL<7708> A_IWL<7707> A_IWL<7706> A_IWL<7705> A_IWL<7704> A_IWL<7703> A_IWL<7702> A_IWL<7701> A_IWL<7700> A_IWL<7699> A_IWL<7698> A_IWL<7697> A_IWL<7696> A_IWL<7695> A_IWL<7694> A_IWL<7693> A_IWL<7692> A_IWL<7691> A_IWL<7690> A_IWL<7689> A_IWL<7688> A_IWL<7687> A_IWL<7686> A_IWL<7685> A_IWL<7684> A_IWL<7683> A_IWL<7682> A_IWL<7681> A_IWL<7680> A_IWL<8191> A_IWL<8190> A_IWL<8189> A_IWL<8188> A_IWL<8187> A_IWL<8186> A_IWL<8185> A_IWL<8184> A_IWL<8183> A_IWL<8182> A_IWL<8181> A_IWL<8180> A_IWL<8179> A_IWL<8178> A_IWL<8177> A_IWL<8176> A_IWL<8175> A_IWL<8174> A_IWL<8173> A_IWL<8172> A_IWL<8171> A_IWL<8170> A_IWL<8169> A_IWL<8168> A_IWL<8167> A_IWL<8166> A_IWL<8165> A_IWL<8164> A_IWL<8163> A_IWL<8162> A_IWL<8161> A_IWL<8160> A_IWL<8159> A_IWL<8158> A_IWL<8157> A_IWL<8156> A_IWL<8155> A_IWL<8154> A_IWL<8153> A_IWL<8152> A_IWL<8151> A_IWL<8150> A_IWL<8149> A_IWL<8148> A_IWL<8147> A_IWL<8146> A_IWL<8145> A_IWL<8144> A_IWL<8143> A_IWL<8142> A_IWL<8141> A_IWL<8140> A_IWL<8139> A_IWL<8138> A_IWL<8137> A_IWL<8136> A_IWL<8135> A_IWL<8134> A_IWL<8133> A_IWL<8132> A_IWL<8131> A_IWL<8130> A_IWL<8129> A_IWL<8128> A_IWL<8127> A_IWL<8126> A_IWL<8125> A_IWL<8124> A_IWL<8123> A_IWL<8122> A_IWL<8121> A_IWL<8120> A_IWL<8119> A_IWL<8118> A_IWL<8117> A_IWL<8116> A_IWL<8115> A_IWL<8114> A_IWL<8113> A_IWL<8112> A_IWL<8111> A_IWL<8110> A_IWL<8109> A_IWL<8108> A_IWL<8107> A_IWL<8106> A_IWL<8105> A_IWL<8104> A_IWL<8103> A_IWL<8102> A_IWL<8101> A_IWL<8100> A_IWL<8099> A_IWL<8098> A_IWL<8097> A_IWL<8096> A_IWL<8095> A_IWL<8094> A_IWL<8093> A_IWL<8092> A_IWL<8091> A_IWL<8090> A_IWL<8089> A_IWL<8088> A_IWL<8087> A_IWL<8086> A_IWL<8085> A_IWL<8084> A_IWL<8083> A_IWL<8082> A_IWL<8081> A_IWL<8080> A_IWL<8079> A_IWL<8078> A_IWL<8077> A_IWL<8076> A_IWL<8075> A_IWL<8074> A_IWL<8073> A_IWL<8072> A_IWL<8071> A_IWL<8070> A_IWL<8069> A_IWL<8068> A_IWL<8067> A_IWL<8066> A_IWL<8065> A_IWL<8064> A_IWL<8063> A_IWL<8062> A_IWL<8061> A_IWL<8060> A_IWL<8059> A_IWL<8058> A_IWL<8057> A_IWL<8056> A_IWL<8055> A_IWL<8054> A_IWL<8053> A_IWL<8052> A_IWL<8051> A_IWL<8050> A_IWL<8049> A_IWL<8048> A_IWL<8047> A_IWL<8046> A_IWL<8045> A_IWL<8044> A_IWL<8043> A_IWL<8042> A_IWL<8041> A_IWL<8040> A_IWL<8039> A_IWL<8038> A_IWL<8037> A_IWL<8036> A_IWL<8035> A_IWL<8034> A_IWL<8033> A_IWL<8032> A_IWL<8031> A_IWL<8030> A_IWL<8029> A_IWL<8028> A_IWL<8027> A_IWL<8026> A_IWL<8025> A_IWL<8024> A_IWL<8023> A_IWL<8022> A_IWL<8021> A_IWL<8020> A_IWL<8019> A_IWL<8018> A_IWL<8017> A_IWL<8016> A_IWL<8015> A_IWL<8014> A_IWL<8013> A_IWL<8012> A_IWL<8011> A_IWL<8010> A_IWL<8009> A_IWL<8008> A_IWL<8007> A_IWL<8006> A_IWL<8005> A_IWL<8004> A_IWL<8003> A_IWL<8002> A_IWL<8001> A_IWL<8000> A_IWL<7999> A_IWL<7998> A_IWL<7997> A_IWL<7996> A_IWL<7995> A_IWL<7994> A_IWL<7993> A_IWL<7992> A_IWL<7991> A_IWL<7990> A_IWL<7989> A_IWL<7988> A_IWL<7987> A_IWL<7986> A_IWL<7985> A_IWL<7984> A_IWL<7983> A_IWL<7982> A_IWL<7981> A_IWL<7980> A_IWL<7979> A_IWL<7978> A_IWL<7977> A_IWL<7976> A_IWL<7975> A_IWL<7974> A_IWL<7973> A_IWL<7972> A_IWL<7971> A_IWL<7970> A_IWL<7969> A_IWL<7968> A_IWL<7967> A_IWL<7966> A_IWL<7965> A_IWL<7964> A_IWL<7963> A_IWL<7962> A_IWL<7961> A_IWL<7960> A_IWL<7959> A_IWL<7958> A_IWL<7957> A_IWL<7956> A_IWL<7955> A_IWL<7954> A_IWL<7953> A_IWL<7952> A_IWL<7951> A_IWL<7950> A_IWL<7949> A_IWL<7948> A_IWL<7947> A_IWL<7946> A_IWL<7945> A_IWL<7944> A_IWL<7943> A_IWL<7942> A_IWL<7941> A_IWL<7940> A_IWL<7939> A_IWL<7938> A_IWL<7937> A_IWL<7936> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<30> A_BLC<61> A_BLC<60> A_BLC_TOP<61> A_BLC_TOP<60> A_BLT<61> A_BLT<60> A_BLT_TOP<61> A_BLT_TOP<60> A_IWL<7679> A_IWL<7678> A_IWL<7677> A_IWL<7676> A_IWL<7675> A_IWL<7674> A_IWL<7673> A_IWL<7672> A_IWL<7671> A_IWL<7670> A_IWL<7669> A_IWL<7668> A_IWL<7667> A_IWL<7666> A_IWL<7665> A_IWL<7664> A_IWL<7663> A_IWL<7662> A_IWL<7661> A_IWL<7660> A_IWL<7659> A_IWL<7658> A_IWL<7657> A_IWL<7656> A_IWL<7655> A_IWL<7654> A_IWL<7653> A_IWL<7652> A_IWL<7651> A_IWL<7650> A_IWL<7649> A_IWL<7648> A_IWL<7647> A_IWL<7646> A_IWL<7645> A_IWL<7644> A_IWL<7643> A_IWL<7642> A_IWL<7641> A_IWL<7640> A_IWL<7639> A_IWL<7638> A_IWL<7637> A_IWL<7636> A_IWL<7635> A_IWL<7634> A_IWL<7633> A_IWL<7632> A_IWL<7631> A_IWL<7630> A_IWL<7629> A_IWL<7628> A_IWL<7627> A_IWL<7626> A_IWL<7625> A_IWL<7624> A_IWL<7623> A_IWL<7622> A_IWL<7621> A_IWL<7620> A_IWL<7619> A_IWL<7618> A_IWL<7617> A_IWL<7616> A_IWL<7615> A_IWL<7614> A_IWL<7613> A_IWL<7612> A_IWL<7611> A_IWL<7610> A_IWL<7609> A_IWL<7608> A_IWL<7607> A_IWL<7606> A_IWL<7605> A_IWL<7604> A_IWL<7603> A_IWL<7602> A_IWL<7601> A_IWL<7600> A_IWL<7599> A_IWL<7598> A_IWL<7597> A_IWL<7596> A_IWL<7595> A_IWL<7594> A_IWL<7593> A_IWL<7592> A_IWL<7591> A_IWL<7590> A_IWL<7589> A_IWL<7588> A_IWL<7587> A_IWL<7586> A_IWL<7585> A_IWL<7584> A_IWL<7583> A_IWL<7582> A_IWL<7581> A_IWL<7580> A_IWL<7579> A_IWL<7578> A_IWL<7577> A_IWL<7576> A_IWL<7575> A_IWL<7574> A_IWL<7573> A_IWL<7572> A_IWL<7571> A_IWL<7570> A_IWL<7569> A_IWL<7568> A_IWL<7567> A_IWL<7566> A_IWL<7565> A_IWL<7564> A_IWL<7563> A_IWL<7562> A_IWL<7561> A_IWL<7560> A_IWL<7559> A_IWL<7558> A_IWL<7557> A_IWL<7556> A_IWL<7555> A_IWL<7554> A_IWL<7553> A_IWL<7552> A_IWL<7551> A_IWL<7550> A_IWL<7549> A_IWL<7548> A_IWL<7547> A_IWL<7546> A_IWL<7545> A_IWL<7544> A_IWL<7543> A_IWL<7542> A_IWL<7541> A_IWL<7540> A_IWL<7539> A_IWL<7538> A_IWL<7537> A_IWL<7536> A_IWL<7535> A_IWL<7534> A_IWL<7533> A_IWL<7532> A_IWL<7531> A_IWL<7530> A_IWL<7529> A_IWL<7528> A_IWL<7527> A_IWL<7526> A_IWL<7525> A_IWL<7524> A_IWL<7523> A_IWL<7522> A_IWL<7521> A_IWL<7520> A_IWL<7519> A_IWL<7518> A_IWL<7517> A_IWL<7516> A_IWL<7515> A_IWL<7514> A_IWL<7513> A_IWL<7512> A_IWL<7511> A_IWL<7510> A_IWL<7509> A_IWL<7508> A_IWL<7507> A_IWL<7506> A_IWL<7505> A_IWL<7504> A_IWL<7503> A_IWL<7502> A_IWL<7501> A_IWL<7500> A_IWL<7499> A_IWL<7498> A_IWL<7497> A_IWL<7496> A_IWL<7495> A_IWL<7494> A_IWL<7493> A_IWL<7492> A_IWL<7491> A_IWL<7490> A_IWL<7489> A_IWL<7488> A_IWL<7487> A_IWL<7486> A_IWL<7485> A_IWL<7484> A_IWL<7483> A_IWL<7482> A_IWL<7481> A_IWL<7480> A_IWL<7479> A_IWL<7478> A_IWL<7477> A_IWL<7476> A_IWL<7475> A_IWL<7474> A_IWL<7473> A_IWL<7472> A_IWL<7471> A_IWL<7470> A_IWL<7469> A_IWL<7468> A_IWL<7467> A_IWL<7466> A_IWL<7465> A_IWL<7464> A_IWL<7463> A_IWL<7462> A_IWL<7461> A_IWL<7460> A_IWL<7459> A_IWL<7458> A_IWL<7457> A_IWL<7456> A_IWL<7455> A_IWL<7454> A_IWL<7453> A_IWL<7452> A_IWL<7451> A_IWL<7450> A_IWL<7449> A_IWL<7448> A_IWL<7447> A_IWL<7446> A_IWL<7445> A_IWL<7444> A_IWL<7443> A_IWL<7442> A_IWL<7441> A_IWL<7440> A_IWL<7439> A_IWL<7438> A_IWL<7437> A_IWL<7436> A_IWL<7435> A_IWL<7434> A_IWL<7433> A_IWL<7432> A_IWL<7431> A_IWL<7430> A_IWL<7429> A_IWL<7428> A_IWL<7427> A_IWL<7426> A_IWL<7425> A_IWL<7424> A_IWL<7935> A_IWL<7934> A_IWL<7933> A_IWL<7932> A_IWL<7931> A_IWL<7930> A_IWL<7929> A_IWL<7928> A_IWL<7927> A_IWL<7926> A_IWL<7925> A_IWL<7924> A_IWL<7923> A_IWL<7922> A_IWL<7921> A_IWL<7920> A_IWL<7919> A_IWL<7918> A_IWL<7917> A_IWL<7916> A_IWL<7915> A_IWL<7914> A_IWL<7913> A_IWL<7912> A_IWL<7911> A_IWL<7910> A_IWL<7909> A_IWL<7908> A_IWL<7907> A_IWL<7906> A_IWL<7905> A_IWL<7904> A_IWL<7903> A_IWL<7902> A_IWL<7901> A_IWL<7900> A_IWL<7899> A_IWL<7898> A_IWL<7897> A_IWL<7896> A_IWL<7895> A_IWL<7894> A_IWL<7893> A_IWL<7892> A_IWL<7891> A_IWL<7890> A_IWL<7889> A_IWL<7888> A_IWL<7887> A_IWL<7886> A_IWL<7885> A_IWL<7884> A_IWL<7883> A_IWL<7882> A_IWL<7881> A_IWL<7880> A_IWL<7879> A_IWL<7878> A_IWL<7877> A_IWL<7876> A_IWL<7875> A_IWL<7874> A_IWL<7873> A_IWL<7872> A_IWL<7871> A_IWL<7870> A_IWL<7869> A_IWL<7868> A_IWL<7867> A_IWL<7866> A_IWL<7865> A_IWL<7864> A_IWL<7863> A_IWL<7862> A_IWL<7861> A_IWL<7860> A_IWL<7859> A_IWL<7858> A_IWL<7857> A_IWL<7856> A_IWL<7855> A_IWL<7854> A_IWL<7853> A_IWL<7852> A_IWL<7851> A_IWL<7850> A_IWL<7849> A_IWL<7848> A_IWL<7847> A_IWL<7846> A_IWL<7845> A_IWL<7844> A_IWL<7843> A_IWL<7842> A_IWL<7841> A_IWL<7840> A_IWL<7839> A_IWL<7838> A_IWL<7837> A_IWL<7836> A_IWL<7835> A_IWL<7834> A_IWL<7833> A_IWL<7832> A_IWL<7831> A_IWL<7830> A_IWL<7829> A_IWL<7828> A_IWL<7827> A_IWL<7826> A_IWL<7825> A_IWL<7824> A_IWL<7823> A_IWL<7822> A_IWL<7821> A_IWL<7820> A_IWL<7819> A_IWL<7818> A_IWL<7817> A_IWL<7816> A_IWL<7815> A_IWL<7814> A_IWL<7813> A_IWL<7812> A_IWL<7811> A_IWL<7810> A_IWL<7809> A_IWL<7808> A_IWL<7807> A_IWL<7806> A_IWL<7805> A_IWL<7804> A_IWL<7803> A_IWL<7802> A_IWL<7801> A_IWL<7800> A_IWL<7799> A_IWL<7798> A_IWL<7797> A_IWL<7796> A_IWL<7795> A_IWL<7794> A_IWL<7793> A_IWL<7792> A_IWL<7791> A_IWL<7790> A_IWL<7789> A_IWL<7788> A_IWL<7787> A_IWL<7786> A_IWL<7785> A_IWL<7784> A_IWL<7783> A_IWL<7782> A_IWL<7781> A_IWL<7780> A_IWL<7779> A_IWL<7778> A_IWL<7777> A_IWL<7776> A_IWL<7775> A_IWL<7774> A_IWL<7773> A_IWL<7772> A_IWL<7771> A_IWL<7770> A_IWL<7769> A_IWL<7768> A_IWL<7767> A_IWL<7766> A_IWL<7765> A_IWL<7764> A_IWL<7763> A_IWL<7762> A_IWL<7761> A_IWL<7760> A_IWL<7759> A_IWL<7758> A_IWL<7757> A_IWL<7756> A_IWL<7755> A_IWL<7754> A_IWL<7753> A_IWL<7752> A_IWL<7751> A_IWL<7750> A_IWL<7749> A_IWL<7748> A_IWL<7747> A_IWL<7746> A_IWL<7745> A_IWL<7744> A_IWL<7743> A_IWL<7742> A_IWL<7741> A_IWL<7740> A_IWL<7739> A_IWL<7738> A_IWL<7737> A_IWL<7736> A_IWL<7735> A_IWL<7734> A_IWL<7733> A_IWL<7732> A_IWL<7731> A_IWL<7730> A_IWL<7729> A_IWL<7728> A_IWL<7727> A_IWL<7726> A_IWL<7725> A_IWL<7724> A_IWL<7723> A_IWL<7722> A_IWL<7721> A_IWL<7720> A_IWL<7719> A_IWL<7718> A_IWL<7717> A_IWL<7716> A_IWL<7715> A_IWL<7714> A_IWL<7713> A_IWL<7712> A_IWL<7711> A_IWL<7710> A_IWL<7709> A_IWL<7708> A_IWL<7707> A_IWL<7706> A_IWL<7705> A_IWL<7704> A_IWL<7703> A_IWL<7702> A_IWL<7701> A_IWL<7700> A_IWL<7699> A_IWL<7698> A_IWL<7697> A_IWL<7696> A_IWL<7695> A_IWL<7694> A_IWL<7693> A_IWL<7692> A_IWL<7691> A_IWL<7690> A_IWL<7689> A_IWL<7688> A_IWL<7687> A_IWL<7686> A_IWL<7685> A_IWL<7684> A_IWL<7683> A_IWL<7682> A_IWL<7681> A_IWL<7680> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<29> A_BLC<59> A_BLC<58> A_BLC_TOP<59> A_BLC_TOP<58> A_BLT<59> A_BLT<58> A_BLT_TOP<59> A_BLT_TOP<58> A_IWL<7423> A_IWL<7422> A_IWL<7421> A_IWL<7420> A_IWL<7419> A_IWL<7418> A_IWL<7417> A_IWL<7416> A_IWL<7415> A_IWL<7414> A_IWL<7413> A_IWL<7412> A_IWL<7411> A_IWL<7410> A_IWL<7409> A_IWL<7408> A_IWL<7407> A_IWL<7406> A_IWL<7405> A_IWL<7404> A_IWL<7403> A_IWL<7402> A_IWL<7401> A_IWL<7400> A_IWL<7399> A_IWL<7398> A_IWL<7397> A_IWL<7396> A_IWL<7395> A_IWL<7394> A_IWL<7393> A_IWL<7392> A_IWL<7391> A_IWL<7390> A_IWL<7389> A_IWL<7388> A_IWL<7387> A_IWL<7386> A_IWL<7385> A_IWL<7384> A_IWL<7383> A_IWL<7382> A_IWL<7381> A_IWL<7380> A_IWL<7379> A_IWL<7378> A_IWL<7377> A_IWL<7376> A_IWL<7375> A_IWL<7374> A_IWL<7373> A_IWL<7372> A_IWL<7371> A_IWL<7370> A_IWL<7369> A_IWL<7368> A_IWL<7367> A_IWL<7366> A_IWL<7365> A_IWL<7364> A_IWL<7363> A_IWL<7362> A_IWL<7361> A_IWL<7360> A_IWL<7359> A_IWL<7358> A_IWL<7357> A_IWL<7356> A_IWL<7355> A_IWL<7354> A_IWL<7353> A_IWL<7352> A_IWL<7351> A_IWL<7350> A_IWL<7349> A_IWL<7348> A_IWL<7347> A_IWL<7346> A_IWL<7345> A_IWL<7344> A_IWL<7343> A_IWL<7342> A_IWL<7341> A_IWL<7340> A_IWL<7339> A_IWL<7338> A_IWL<7337> A_IWL<7336> A_IWL<7335> A_IWL<7334> A_IWL<7333> A_IWL<7332> A_IWL<7331> A_IWL<7330> A_IWL<7329> A_IWL<7328> A_IWL<7327> A_IWL<7326> A_IWL<7325> A_IWL<7324> A_IWL<7323> A_IWL<7322> A_IWL<7321> A_IWL<7320> A_IWL<7319> A_IWL<7318> A_IWL<7317> A_IWL<7316> A_IWL<7315> A_IWL<7314> A_IWL<7313> A_IWL<7312> A_IWL<7311> A_IWL<7310> A_IWL<7309> A_IWL<7308> A_IWL<7307> A_IWL<7306> A_IWL<7305> A_IWL<7304> A_IWL<7303> A_IWL<7302> A_IWL<7301> A_IWL<7300> A_IWL<7299> A_IWL<7298> A_IWL<7297> A_IWL<7296> A_IWL<7295> A_IWL<7294> A_IWL<7293> A_IWL<7292> A_IWL<7291> A_IWL<7290> A_IWL<7289> A_IWL<7288> A_IWL<7287> A_IWL<7286> A_IWL<7285> A_IWL<7284> A_IWL<7283> A_IWL<7282> A_IWL<7281> A_IWL<7280> A_IWL<7279> A_IWL<7278> A_IWL<7277> A_IWL<7276> A_IWL<7275> A_IWL<7274> A_IWL<7273> A_IWL<7272> A_IWL<7271> A_IWL<7270> A_IWL<7269> A_IWL<7268> A_IWL<7267> A_IWL<7266> A_IWL<7265> A_IWL<7264> A_IWL<7263> A_IWL<7262> A_IWL<7261> A_IWL<7260> A_IWL<7259> A_IWL<7258> A_IWL<7257> A_IWL<7256> A_IWL<7255> A_IWL<7254> A_IWL<7253> A_IWL<7252> A_IWL<7251> A_IWL<7250> A_IWL<7249> A_IWL<7248> A_IWL<7247> A_IWL<7246> A_IWL<7245> A_IWL<7244> A_IWL<7243> A_IWL<7242> A_IWL<7241> A_IWL<7240> A_IWL<7239> A_IWL<7238> A_IWL<7237> A_IWL<7236> A_IWL<7235> A_IWL<7234> A_IWL<7233> A_IWL<7232> A_IWL<7231> A_IWL<7230> A_IWL<7229> A_IWL<7228> A_IWL<7227> A_IWL<7226> A_IWL<7225> A_IWL<7224> A_IWL<7223> A_IWL<7222> A_IWL<7221> A_IWL<7220> A_IWL<7219> A_IWL<7218> A_IWL<7217> A_IWL<7216> A_IWL<7215> A_IWL<7214> A_IWL<7213> A_IWL<7212> A_IWL<7211> A_IWL<7210> A_IWL<7209> A_IWL<7208> A_IWL<7207> A_IWL<7206> A_IWL<7205> A_IWL<7204> A_IWL<7203> A_IWL<7202> A_IWL<7201> A_IWL<7200> A_IWL<7199> A_IWL<7198> A_IWL<7197> A_IWL<7196> A_IWL<7195> A_IWL<7194> A_IWL<7193> A_IWL<7192> A_IWL<7191> A_IWL<7190> A_IWL<7189> A_IWL<7188> A_IWL<7187> A_IWL<7186> A_IWL<7185> A_IWL<7184> A_IWL<7183> A_IWL<7182> A_IWL<7181> A_IWL<7180> A_IWL<7179> A_IWL<7178> A_IWL<7177> A_IWL<7176> A_IWL<7175> A_IWL<7174> A_IWL<7173> A_IWL<7172> A_IWL<7171> A_IWL<7170> A_IWL<7169> A_IWL<7168> A_IWL<7679> A_IWL<7678> A_IWL<7677> A_IWL<7676> A_IWL<7675> A_IWL<7674> A_IWL<7673> A_IWL<7672> A_IWL<7671> A_IWL<7670> A_IWL<7669> A_IWL<7668> A_IWL<7667> A_IWL<7666> A_IWL<7665> A_IWL<7664> A_IWL<7663> A_IWL<7662> A_IWL<7661> A_IWL<7660> A_IWL<7659> A_IWL<7658> A_IWL<7657> A_IWL<7656> A_IWL<7655> A_IWL<7654> A_IWL<7653> A_IWL<7652> A_IWL<7651> A_IWL<7650> A_IWL<7649> A_IWL<7648> A_IWL<7647> A_IWL<7646> A_IWL<7645> A_IWL<7644> A_IWL<7643> A_IWL<7642> A_IWL<7641> A_IWL<7640> A_IWL<7639> A_IWL<7638> A_IWL<7637> A_IWL<7636> A_IWL<7635> A_IWL<7634> A_IWL<7633> A_IWL<7632> A_IWL<7631> A_IWL<7630> A_IWL<7629> A_IWL<7628> A_IWL<7627> A_IWL<7626> A_IWL<7625> A_IWL<7624> A_IWL<7623> A_IWL<7622> A_IWL<7621> A_IWL<7620> A_IWL<7619> A_IWL<7618> A_IWL<7617> A_IWL<7616> A_IWL<7615> A_IWL<7614> A_IWL<7613> A_IWL<7612> A_IWL<7611> A_IWL<7610> A_IWL<7609> A_IWL<7608> A_IWL<7607> A_IWL<7606> A_IWL<7605> A_IWL<7604> A_IWL<7603> A_IWL<7602> A_IWL<7601> A_IWL<7600> A_IWL<7599> A_IWL<7598> A_IWL<7597> A_IWL<7596> A_IWL<7595> A_IWL<7594> A_IWL<7593> A_IWL<7592> A_IWL<7591> A_IWL<7590> A_IWL<7589> A_IWL<7588> A_IWL<7587> A_IWL<7586> A_IWL<7585> A_IWL<7584> A_IWL<7583> A_IWL<7582> A_IWL<7581> A_IWL<7580> A_IWL<7579> A_IWL<7578> A_IWL<7577> A_IWL<7576> A_IWL<7575> A_IWL<7574> A_IWL<7573> A_IWL<7572> A_IWL<7571> A_IWL<7570> A_IWL<7569> A_IWL<7568> A_IWL<7567> A_IWL<7566> A_IWL<7565> A_IWL<7564> A_IWL<7563> A_IWL<7562> A_IWL<7561> A_IWL<7560> A_IWL<7559> A_IWL<7558> A_IWL<7557> A_IWL<7556> A_IWL<7555> A_IWL<7554> A_IWL<7553> A_IWL<7552> A_IWL<7551> A_IWL<7550> A_IWL<7549> A_IWL<7548> A_IWL<7547> A_IWL<7546> A_IWL<7545> A_IWL<7544> A_IWL<7543> A_IWL<7542> A_IWL<7541> A_IWL<7540> A_IWL<7539> A_IWL<7538> A_IWL<7537> A_IWL<7536> A_IWL<7535> A_IWL<7534> A_IWL<7533> A_IWL<7532> A_IWL<7531> A_IWL<7530> A_IWL<7529> A_IWL<7528> A_IWL<7527> A_IWL<7526> A_IWL<7525> A_IWL<7524> A_IWL<7523> A_IWL<7522> A_IWL<7521> A_IWL<7520> A_IWL<7519> A_IWL<7518> A_IWL<7517> A_IWL<7516> A_IWL<7515> A_IWL<7514> A_IWL<7513> A_IWL<7512> A_IWL<7511> A_IWL<7510> A_IWL<7509> A_IWL<7508> A_IWL<7507> A_IWL<7506> A_IWL<7505> A_IWL<7504> A_IWL<7503> A_IWL<7502> A_IWL<7501> A_IWL<7500> A_IWL<7499> A_IWL<7498> A_IWL<7497> A_IWL<7496> A_IWL<7495> A_IWL<7494> A_IWL<7493> A_IWL<7492> A_IWL<7491> A_IWL<7490> A_IWL<7489> A_IWL<7488> A_IWL<7487> A_IWL<7486> A_IWL<7485> A_IWL<7484> A_IWL<7483> A_IWL<7482> A_IWL<7481> A_IWL<7480> A_IWL<7479> A_IWL<7478> A_IWL<7477> A_IWL<7476> A_IWL<7475> A_IWL<7474> A_IWL<7473> A_IWL<7472> A_IWL<7471> A_IWL<7470> A_IWL<7469> A_IWL<7468> A_IWL<7467> A_IWL<7466> A_IWL<7465> A_IWL<7464> A_IWL<7463> A_IWL<7462> A_IWL<7461> A_IWL<7460> A_IWL<7459> A_IWL<7458> A_IWL<7457> A_IWL<7456> A_IWL<7455> A_IWL<7454> A_IWL<7453> A_IWL<7452> A_IWL<7451> A_IWL<7450> A_IWL<7449> A_IWL<7448> A_IWL<7447> A_IWL<7446> A_IWL<7445> A_IWL<7444> A_IWL<7443> A_IWL<7442> A_IWL<7441> A_IWL<7440> A_IWL<7439> A_IWL<7438> A_IWL<7437> A_IWL<7436> A_IWL<7435> A_IWL<7434> A_IWL<7433> A_IWL<7432> A_IWL<7431> A_IWL<7430> A_IWL<7429> A_IWL<7428> A_IWL<7427> A_IWL<7426> A_IWL<7425> A_IWL<7424> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<28> A_BLC<57> A_BLC<56> A_BLC_TOP<57> A_BLC_TOP<56> A_BLT<57> A_BLT<56> A_BLT_TOP<57> A_BLT_TOP<56> A_IWL<7167> A_IWL<7166> A_IWL<7165> A_IWL<7164> A_IWL<7163> A_IWL<7162> A_IWL<7161> A_IWL<7160> A_IWL<7159> A_IWL<7158> A_IWL<7157> A_IWL<7156> A_IWL<7155> A_IWL<7154> A_IWL<7153> A_IWL<7152> A_IWL<7151> A_IWL<7150> A_IWL<7149> A_IWL<7148> A_IWL<7147> A_IWL<7146> A_IWL<7145> A_IWL<7144> A_IWL<7143> A_IWL<7142> A_IWL<7141> A_IWL<7140> A_IWL<7139> A_IWL<7138> A_IWL<7137> A_IWL<7136> A_IWL<7135> A_IWL<7134> A_IWL<7133> A_IWL<7132> A_IWL<7131> A_IWL<7130> A_IWL<7129> A_IWL<7128> A_IWL<7127> A_IWL<7126> A_IWL<7125> A_IWL<7124> A_IWL<7123> A_IWL<7122> A_IWL<7121> A_IWL<7120> A_IWL<7119> A_IWL<7118> A_IWL<7117> A_IWL<7116> A_IWL<7115> A_IWL<7114> A_IWL<7113> A_IWL<7112> A_IWL<7111> A_IWL<7110> A_IWL<7109> A_IWL<7108> A_IWL<7107> A_IWL<7106> A_IWL<7105> A_IWL<7104> A_IWL<7103> A_IWL<7102> A_IWL<7101> A_IWL<7100> A_IWL<7099> A_IWL<7098> A_IWL<7097> A_IWL<7096> A_IWL<7095> A_IWL<7094> A_IWL<7093> A_IWL<7092> A_IWL<7091> A_IWL<7090> A_IWL<7089> A_IWL<7088> A_IWL<7087> A_IWL<7086> A_IWL<7085> A_IWL<7084> A_IWL<7083> A_IWL<7082> A_IWL<7081> A_IWL<7080> A_IWL<7079> A_IWL<7078> A_IWL<7077> A_IWL<7076> A_IWL<7075> A_IWL<7074> A_IWL<7073> A_IWL<7072> A_IWL<7071> A_IWL<7070> A_IWL<7069> A_IWL<7068> A_IWL<7067> A_IWL<7066> A_IWL<7065> A_IWL<7064> A_IWL<7063> A_IWL<7062> A_IWL<7061> A_IWL<7060> A_IWL<7059> A_IWL<7058> A_IWL<7057> A_IWL<7056> A_IWL<7055> A_IWL<7054> A_IWL<7053> A_IWL<7052> A_IWL<7051> A_IWL<7050> A_IWL<7049> A_IWL<7048> A_IWL<7047> A_IWL<7046> A_IWL<7045> A_IWL<7044> A_IWL<7043> A_IWL<7042> A_IWL<7041> A_IWL<7040> A_IWL<7039> A_IWL<7038> A_IWL<7037> A_IWL<7036> A_IWL<7035> A_IWL<7034> A_IWL<7033> A_IWL<7032> A_IWL<7031> A_IWL<7030> A_IWL<7029> A_IWL<7028> A_IWL<7027> A_IWL<7026> A_IWL<7025> A_IWL<7024> A_IWL<7023> A_IWL<7022> A_IWL<7021> A_IWL<7020> A_IWL<7019> A_IWL<7018> A_IWL<7017> A_IWL<7016> A_IWL<7015> A_IWL<7014> A_IWL<7013> A_IWL<7012> A_IWL<7011> A_IWL<7010> A_IWL<7009> A_IWL<7008> A_IWL<7007> A_IWL<7006> A_IWL<7005> A_IWL<7004> A_IWL<7003> A_IWL<7002> A_IWL<7001> A_IWL<7000> A_IWL<6999> A_IWL<6998> A_IWL<6997> A_IWL<6996> A_IWL<6995> A_IWL<6994> A_IWL<6993> A_IWL<6992> A_IWL<6991> A_IWL<6990> A_IWL<6989> A_IWL<6988> A_IWL<6987> A_IWL<6986> A_IWL<6985> A_IWL<6984> A_IWL<6983> A_IWL<6982> A_IWL<6981> A_IWL<6980> A_IWL<6979> A_IWL<6978> A_IWL<6977> A_IWL<6976> A_IWL<6975> A_IWL<6974> A_IWL<6973> A_IWL<6972> A_IWL<6971> A_IWL<6970> A_IWL<6969> A_IWL<6968> A_IWL<6967> A_IWL<6966> A_IWL<6965> A_IWL<6964> A_IWL<6963> A_IWL<6962> A_IWL<6961> A_IWL<6960> A_IWL<6959> A_IWL<6958> A_IWL<6957> A_IWL<6956> A_IWL<6955> A_IWL<6954> A_IWL<6953> A_IWL<6952> A_IWL<6951> A_IWL<6950> A_IWL<6949> A_IWL<6948> A_IWL<6947> A_IWL<6946> A_IWL<6945> A_IWL<6944> A_IWL<6943> A_IWL<6942> A_IWL<6941> A_IWL<6940> A_IWL<6939> A_IWL<6938> A_IWL<6937> A_IWL<6936> A_IWL<6935> A_IWL<6934> A_IWL<6933> A_IWL<6932> A_IWL<6931> A_IWL<6930> A_IWL<6929> A_IWL<6928> A_IWL<6927> A_IWL<6926> A_IWL<6925> A_IWL<6924> A_IWL<6923> A_IWL<6922> A_IWL<6921> A_IWL<6920> A_IWL<6919> A_IWL<6918> A_IWL<6917> A_IWL<6916> A_IWL<6915> A_IWL<6914> A_IWL<6913> A_IWL<6912> A_IWL<7423> A_IWL<7422> A_IWL<7421> A_IWL<7420> A_IWL<7419> A_IWL<7418> A_IWL<7417> A_IWL<7416> A_IWL<7415> A_IWL<7414> A_IWL<7413> A_IWL<7412> A_IWL<7411> A_IWL<7410> A_IWL<7409> A_IWL<7408> A_IWL<7407> A_IWL<7406> A_IWL<7405> A_IWL<7404> A_IWL<7403> A_IWL<7402> A_IWL<7401> A_IWL<7400> A_IWL<7399> A_IWL<7398> A_IWL<7397> A_IWL<7396> A_IWL<7395> A_IWL<7394> A_IWL<7393> A_IWL<7392> A_IWL<7391> A_IWL<7390> A_IWL<7389> A_IWL<7388> A_IWL<7387> A_IWL<7386> A_IWL<7385> A_IWL<7384> A_IWL<7383> A_IWL<7382> A_IWL<7381> A_IWL<7380> A_IWL<7379> A_IWL<7378> A_IWL<7377> A_IWL<7376> A_IWL<7375> A_IWL<7374> A_IWL<7373> A_IWL<7372> A_IWL<7371> A_IWL<7370> A_IWL<7369> A_IWL<7368> A_IWL<7367> A_IWL<7366> A_IWL<7365> A_IWL<7364> A_IWL<7363> A_IWL<7362> A_IWL<7361> A_IWL<7360> A_IWL<7359> A_IWL<7358> A_IWL<7357> A_IWL<7356> A_IWL<7355> A_IWL<7354> A_IWL<7353> A_IWL<7352> A_IWL<7351> A_IWL<7350> A_IWL<7349> A_IWL<7348> A_IWL<7347> A_IWL<7346> A_IWL<7345> A_IWL<7344> A_IWL<7343> A_IWL<7342> A_IWL<7341> A_IWL<7340> A_IWL<7339> A_IWL<7338> A_IWL<7337> A_IWL<7336> A_IWL<7335> A_IWL<7334> A_IWL<7333> A_IWL<7332> A_IWL<7331> A_IWL<7330> A_IWL<7329> A_IWL<7328> A_IWL<7327> A_IWL<7326> A_IWL<7325> A_IWL<7324> A_IWL<7323> A_IWL<7322> A_IWL<7321> A_IWL<7320> A_IWL<7319> A_IWL<7318> A_IWL<7317> A_IWL<7316> A_IWL<7315> A_IWL<7314> A_IWL<7313> A_IWL<7312> A_IWL<7311> A_IWL<7310> A_IWL<7309> A_IWL<7308> A_IWL<7307> A_IWL<7306> A_IWL<7305> A_IWL<7304> A_IWL<7303> A_IWL<7302> A_IWL<7301> A_IWL<7300> A_IWL<7299> A_IWL<7298> A_IWL<7297> A_IWL<7296> A_IWL<7295> A_IWL<7294> A_IWL<7293> A_IWL<7292> A_IWL<7291> A_IWL<7290> A_IWL<7289> A_IWL<7288> A_IWL<7287> A_IWL<7286> A_IWL<7285> A_IWL<7284> A_IWL<7283> A_IWL<7282> A_IWL<7281> A_IWL<7280> A_IWL<7279> A_IWL<7278> A_IWL<7277> A_IWL<7276> A_IWL<7275> A_IWL<7274> A_IWL<7273> A_IWL<7272> A_IWL<7271> A_IWL<7270> A_IWL<7269> A_IWL<7268> A_IWL<7267> A_IWL<7266> A_IWL<7265> A_IWL<7264> A_IWL<7263> A_IWL<7262> A_IWL<7261> A_IWL<7260> A_IWL<7259> A_IWL<7258> A_IWL<7257> A_IWL<7256> A_IWL<7255> A_IWL<7254> A_IWL<7253> A_IWL<7252> A_IWL<7251> A_IWL<7250> A_IWL<7249> A_IWL<7248> A_IWL<7247> A_IWL<7246> A_IWL<7245> A_IWL<7244> A_IWL<7243> A_IWL<7242> A_IWL<7241> A_IWL<7240> A_IWL<7239> A_IWL<7238> A_IWL<7237> A_IWL<7236> A_IWL<7235> A_IWL<7234> A_IWL<7233> A_IWL<7232> A_IWL<7231> A_IWL<7230> A_IWL<7229> A_IWL<7228> A_IWL<7227> A_IWL<7226> A_IWL<7225> A_IWL<7224> A_IWL<7223> A_IWL<7222> A_IWL<7221> A_IWL<7220> A_IWL<7219> A_IWL<7218> A_IWL<7217> A_IWL<7216> A_IWL<7215> A_IWL<7214> A_IWL<7213> A_IWL<7212> A_IWL<7211> A_IWL<7210> A_IWL<7209> A_IWL<7208> A_IWL<7207> A_IWL<7206> A_IWL<7205> A_IWL<7204> A_IWL<7203> A_IWL<7202> A_IWL<7201> A_IWL<7200> A_IWL<7199> A_IWL<7198> A_IWL<7197> A_IWL<7196> A_IWL<7195> A_IWL<7194> A_IWL<7193> A_IWL<7192> A_IWL<7191> A_IWL<7190> A_IWL<7189> A_IWL<7188> A_IWL<7187> A_IWL<7186> A_IWL<7185> A_IWL<7184> A_IWL<7183> A_IWL<7182> A_IWL<7181> A_IWL<7180> A_IWL<7179> A_IWL<7178> A_IWL<7177> A_IWL<7176> A_IWL<7175> A_IWL<7174> A_IWL<7173> A_IWL<7172> A_IWL<7171> A_IWL<7170> A_IWL<7169> A_IWL<7168> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<27> A_BLC<55> A_BLC<54> A_BLC_TOP<55> A_BLC_TOP<54> A_BLT<55> A_BLT<54> A_BLT_TOP<55> A_BLT_TOP<54> A_IWL<6911> A_IWL<6910> A_IWL<6909> A_IWL<6908> A_IWL<6907> A_IWL<6906> A_IWL<6905> A_IWL<6904> A_IWL<6903> A_IWL<6902> A_IWL<6901> A_IWL<6900> A_IWL<6899> A_IWL<6898> A_IWL<6897> A_IWL<6896> A_IWL<6895> A_IWL<6894> A_IWL<6893> A_IWL<6892> A_IWL<6891> A_IWL<6890> A_IWL<6889> A_IWL<6888> A_IWL<6887> A_IWL<6886> A_IWL<6885> A_IWL<6884> A_IWL<6883> A_IWL<6882> A_IWL<6881> A_IWL<6880> A_IWL<6879> A_IWL<6878> A_IWL<6877> A_IWL<6876> A_IWL<6875> A_IWL<6874> A_IWL<6873> A_IWL<6872> A_IWL<6871> A_IWL<6870> A_IWL<6869> A_IWL<6868> A_IWL<6867> A_IWL<6866> A_IWL<6865> A_IWL<6864> A_IWL<6863> A_IWL<6862> A_IWL<6861> A_IWL<6860> A_IWL<6859> A_IWL<6858> A_IWL<6857> A_IWL<6856> A_IWL<6855> A_IWL<6854> A_IWL<6853> A_IWL<6852> A_IWL<6851> A_IWL<6850> A_IWL<6849> A_IWL<6848> A_IWL<6847> A_IWL<6846> A_IWL<6845> A_IWL<6844> A_IWL<6843> A_IWL<6842> A_IWL<6841> A_IWL<6840> A_IWL<6839> A_IWL<6838> A_IWL<6837> A_IWL<6836> A_IWL<6835> A_IWL<6834> A_IWL<6833> A_IWL<6832> A_IWL<6831> A_IWL<6830> A_IWL<6829> A_IWL<6828> A_IWL<6827> A_IWL<6826> A_IWL<6825> A_IWL<6824> A_IWL<6823> A_IWL<6822> A_IWL<6821> A_IWL<6820> A_IWL<6819> A_IWL<6818> A_IWL<6817> A_IWL<6816> A_IWL<6815> A_IWL<6814> A_IWL<6813> A_IWL<6812> A_IWL<6811> A_IWL<6810> A_IWL<6809> A_IWL<6808> A_IWL<6807> A_IWL<6806> A_IWL<6805> A_IWL<6804> A_IWL<6803> A_IWL<6802> A_IWL<6801> A_IWL<6800> A_IWL<6799> A_IWL<6798> A_IWL<6797> A_IWL<6796> A_IWL<6795> A_IWL<6794> A_IWL<6793> A_IWL<6792> A_IWL<6791> A_IWL<6790> A_IWL<6789> A_IWL<6788> A_IWL<6787> A_IWL<6786> A_IWL<6785> A_IWL<6784> A_IWL<6783> A_IWL<6782> A_IWL<6781> A_IWL<6780> A_IWL<6779> A_IWL<6778> A_IWL<6777> A_IWL<6776> A_IWL<6775> A_IWL<6774> A_IWL<6773> A_IWL<6772> A_IWL<6771> A_IWL<6770> A_IWL<6769> A_IWL<6768> A_IWL<6767> A_IWL<6766> A_IWL<6765> A_IWL<6764> A_IWL<6763> A_IWL<6762> A_IWL<6761> A_IWL<6760> A_IWL<6759> A_IWL<6758> A_IWL<6757> A_IWL<6756> A_IWL<6755> A_IWL<6754> A_IWL<6753> A_IWL<6752> A_IWL<6751> A_IWL<6750> A_IWL<6749> A_IWL<6748> A_IWL<6747> A_IWL<6746> A_IWL<6745> A_IWL<6744> A_IWL<6743> A_IWL<6742> A_IWL<6741> A_IWL<6740> A_IWL<6739> A_IWL<6738> A_IWL<6737> A_IWL<6736> A_IWL<6735> A_IWL<6734> A_IWL<6733> A_IWL<6732> A_IWL<6731> A_IWL<6730> A_IWL<6729> A_IWL<6728> A_IWL<6727> A_IWL<6726> A_IWL<6725> A_IWL<6724> A_IWL<6723> A_IWL<6722> A_IWL<6721> A_IWL<6720> A_IWL<6719> A_IWL<6718> A_IWL<6717> A_IWL<6716> A_IWL<6715> A_IWL<6714> A_IWL<6713> A_IWL<6712> A_IWL<6711> A_IWL<6710> A_IWL<6709> A_IWL<6708> A_IWL<6707> A_IWL<6706> A_IWL<6705> A_IWL<6704> A_IWL<6703> A_IWL<6702> A_IWL<6701> A_IWL<6700> A_IWL<6699> A_IWL<6698> A_IWL<6697> A_IWL<6696> A_IWL<6695> A_IWL<6694> A_IWL<6693> A_IWL<6692> A_IWL<6691> A_IWL<6690> A_IWL<6689> A_IWL<6688> A_IWL<6687> A_IWL<6686> A_IWL<6685> A_IWL<6684> A_IWL<6683> A_IWL<6682> A_IWL<6681> A_IWL<6680> A_IWL<6679> A_IWL<6678> A_IWL<6677> A_IWL<6676> A_IWL<6675> A_IWL<6674> A_IWL<6673> A_IWL<6672> A_IWL<6671> A_IWL<6670> A_IWL<6669> A_IWL<6668> A_IWL<6667> A_IWL<6666> A_IWL<6665> A_IWL<6664> A_IWL<6663> A_IWL<6662> A_IWL<6661> A_IWL<6660> A_IWL<6659> A_IWL<6658> A_IWL<6657> A_IWL<6656> A_IWL<7167> A_IWL<7166> A_IWL<7165> A_IWL<7164> A_IWL<7163> A_IWL<7162> A_IWL<7161> A_IWL<7160> A_IWL<7159> A_IWL<7158> A_IWL<7157> A_IWL<7156> A_IWL<7155> A_IWL<7154> A_IWL<7153> A_IWL<7152> A_IWL<7151> A_IWL<7150> A_IWL<7149> A_IWL<7148> A_IWL<7147> A_IWL<7146> A_IWL<7145> A_IWL<7144> A_IWL<7143> A_IWL<7142> A_IWL<7141> A_IWL<7140> A_IWL<7139> A_IWL<7138> A_IWL<7137> A_IWL<7136> A_IWL<7135> A_IWL<7134> A_IWL<7133> A_IWL<7132> A_IWL<7131> A_IWL<7130> A_IWL<7129> A_IWL<7128> A_IWL<7127> A_IWL<7126> A_IWL<7125> A_IWL<7124> A_IWL<7123> A_IWL<7122> A_IWL<7121> A_IWL<7120> A_IWL<7119> A_IWL<7118> A_IWL<7117> A_IWL<7116> A_IWL<7115> A_IWL<7114> A_IWL<7113> A_IWL<7112> A_IWL<7111> A_IWL<7110> A_IWL<7109> A_IWL<7108> A_IWL<7107> A_IWL<7106> A_IWL<7105> A_IWL<7104> A_IWL<7103> A_IWL<7102> A_IWL<7101> A_IWL<7100> A_IWL<7099> A_IWL<7098> A_IWL<7097> A_IWL<7096> A_IWL<7095> A_IWL<7094> A_IWL<7093> A_IWL<7092> A_IWL<7091> A_IWL<7090> A_IWL<7089> A_IWL<7088> A_IWL<7087> A_IWL<7086> A_IWL<7085> A_IWL<7084> A_IWL<7083> A_IWL<7082> A_IWL<7081> A_IWL<7080> A_IWL<7079> A_IWL<7078> A_IWL<7077> A_IWL<7076> A_IWL<7075> A_IWL<7074> A_IWL<7073> A_IWL<7072> A_IWL<7071> A_IWL<7070> A_IWL<7069> A_IWL<7068> A_IWL<7067> A_IWL<7066> A_IWL<7065> A_IWL<7064> A_IWL<7063> A_IWL<7062> A_IWL<7061> A_IWL<7060> A_IWL<7059> A_IWL<7058> A_IWL<7057> A_IWL<7056> A_IWL<7055> A_IWL<7054> A_IWL<7053> A_IWL<7052> A_IWL<7051> A_IWL<7050> A_IWL<7049> A_IWL<7048> A_IWL<7047> A_IWL<7046> A_IWL<7045> A_IWL<7044> A_IWL<7043> A_IWL<7042> A_IWL<7041> A_IWL<7040> A_IWL<7039> A_IWL<7038> A_IWL<7037> A_IWL<7036> A_IWL<7035> A_IWL<7034> A_IWL<7033> A_IWL<7032> A_IWL<7031> A_IWL<7030> A_IWL<7029> A_IWL<7028> A_IWL<7027> A_IWL<7026> A_IWL<7025> A_IWL<7024> A_IWL<7023> A_IWL<7022> A_IWL<7021> A_IWL<7020> A_IWL<7019> A_IWL<7018> A_IWL<7017> A_IWL<7016> A_IWL<7015> A_IWL<7014> A_IWL<7013> A_IWL<7012> A_IWL<7011> A_IWL<7010> A_IWL<7009> A_IWL<7008> A_IWL<7007> A_IWL<7006> A_IWL<7005> A_IWL<7004> A_IWL<7003> A_IWL<7002> A_IWL<7001> A_IWL<7000> A_IWL<6999> A_IWL<6998> A_IWL<6997> A_IWL<6996> A_IWL<6995> A_IWL<6994> A_IWL<6993> A_IWL<6992> A_IWL<6991> A_IWL<6990> A_IWL<6989> A_IWL<6988> A_IWL<6987> A_IWL<6986> A_IWL<6985> A_IWL<6984> A_IWL<6983> A_IWL<6982> A_IWL<6981> A_IWL<6980> A_IWL<6979> A_IWL<6978> A_IWL<6977> A_IWL<6976> A_IWL<6975> A_IWL<6974> A_IWL<6973> A_IWL<6972> A_IWL<6971> A_IWL<6970> A_IWL<6969> A_IWL<6968> A_IWL<6967> A_IWL<6966> A_IWL<6965> A_IWL<6964> A_IWL<6963> A_IWL<6962> A_IWL<6961> A_IWL<6960> A_IWL<6959> A_IWL<6958> A_IWL<6957> A_IWL<6956> A_IWL<6955> A_IWL<6954> A_IWL<6953> A_IWL<6952> A_IWL<6951> A_IWL<6950> A_IWL<6949> A_IWL<6948> A_IWL<6947> A_IWL<6946> A_IWL<6945> A_IWL<6944> A_IWL<6943> A_IWL<6942> A_IWL<6941> A_IWL<6940> A_IWL<6939> A_IWL<6938> A_IWL<6937> A_IWL<6936> A_IWL<6935> A_IWL<6934> A_IWL<6933> A_IWL<6932> A_IWL<6931> A_IWL<6930> A_IWL<6929> A_IWL<6928> A_IWL<6927> A_IWL<6926> A_IWL<6925> A_IWL<6924> A_IWL<6923> A_IWL<6922> A_IWL<6921> A_IWL<6920> A_IWL<6919> A_IWL<6918> A_IWL<6917> A_IWL<6916> A_IWL<6915> A_IWL<6914> A_IWL<6913> A_IWL<6912> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<26> A_BLC<53> A_BLC<52> A_BLC_TOP<53> A_BLC_TOP<52> A_BLT<53> A_BLT<52> A_BLT_TOP<53> A_BLT_TOP<52> A_IWL<6655> A_IWL<6654> A_IWL<6653> A_IWL<6652> A_IWL<6651> A_IWL<6650> A_IWL<6649> A_IWL<6648> A_IWL<6647> A_IWL<6646> A_IWL<6645> A_IWL<6644> A_IWL<6643> A_IWL<6642> A_IWL<6641> A_IWL<6640> A_IWL<6639> A_IWL<6638> A_IWL<6637> A_IWL<6636> A_IWL<6635> A_IWL<6634> A_IWL<6633> A_IWL<6632> A_IWL<6631> A_IWL<6630> A_IWL<6629> A_IWL<6628> A_IWL<6627> A_IWL<6626> A_IWL<6625> A_IWL<6624> A_IWL<6623> A_IWL<6622> A_IWL<6621> A_IWL<6620> A_IWL<6619> A_IWL<6618> A_IWL<6617> A_IWL<6616> A_IWL<6615> A_IWL<6614> A_IWL<6613> A_IWL<6612> A_IWL<6611> A_IWL<6610> A_IWL<6609> A_IWL<6608> A_IWL<6607> A_IWL<6606> A_IWL<6605> A_IWL<6604> A_IWL<6603> A_IWL<6602> A_IWL<6601> A_IWL<6600> A_IWL<6599> A_IWL<6598> A_IWL<6597> A_IWL<6596> A_IWL<6595> A_IWL<6594> A_IWL<6593> A_IWL<6592> A_IWL<6591> A_IWL<6590> A_IWL<6589> A_IWL<6588> A_IWL<6587> A_IWL<6586> A_IWL<6585> A_IWL<6584> A_IWL<6583> A_IWL<6582> A_IWL<6581> A_IWL<6580> A_IWL<6579> A_IWL<6578> A_IWL<6577> A_IWL<6576> A_IWL<6575> A_IWL<6574> A_IWL<6573> A_IWL<6572> A_IWL<6571> A_IWL<6570> A_IWL<6569> A_IWL<6568> A_IWL<6567> A_IWL<6566> A_IWL<6565> A_IWL<6564> A_IWL<6563> A_IWL<6562> A_IWL<6561> A_IWL<6560> A_IWL<6559> A_IWL<6558> A_IWL<6557> A_IWL<6556> A_IWL<6555> A_IWL<6554> A_IWL<6553> A_IWL<6552> A_IWL<6551> A_IWL<6550> A_IWL<6549> A_IWL<6548> A_IWL<6547> A_IWL<6546> A_IWL<6545> A_IWL<6544> A_IWL<6543> A_IWL<6542> A_IWL<6541> A_IWL<6540> A_IWL<6539> A_IWL<6538> A_IWL<6537> A_IWL<6536> A_IWL<6535> A_IWL<6534> A_IWL<6533> A_IWL<6532> A_IWL<6531> A_IWL<6530> A_IWL<6529> A_IWL<6528> A_IWL<6527> A_IWL<6526> A_IWL<6525> A_IWL<6524> A_IWL<6523> A_IWL<6522> A_IWL<6521> A_IWL<6520> A_IWL<6519> A_IWL<6518> A_IWL<6517> A_IWL<6516> A_IWL<6515> A_IWL<6514> A_IWL<6513> A_IWL<6512> A_IWL<6511> A_IWL<6510> A_IWL<6509> A_IWL<6508> A_IWL<6507> A_IWL<6506> A_IWL<6505> A_IWL<6504> A_IWL<6503> A_IWL<6502> A_IWL<6501> A_IWL<6500> A_IWL<6499> A_IWL<6498> A_IWL<6497> A_IWL<6496> A_IWL<6495> A_IWL<6494> A_IWL<6493> A_IWL<6492> A_IWL<6491> A_IWL<6490> A_IWL<6489> A_IWL<6488> A_IWL<6487> A_IWL<6486> A_IWL<6485> A_IWL<6484> A_IWL<6483> A_IWL<6482> A_IWL<6481> A_IWL<6480> A_IWL<6479> A_IWL<6478> A_IWL<6477> A_IWL<6476> A_IWL<6475> A_IWL<6474> A_IWL<6473> A_IWL<6472> A_IWL<6471> A_IWL<6470> A_IWL<6469> A_IWL<6468> A_IWL<6467> A_IWL<6466> A_IWL<6465> A_IWL<6464> A_IWL<6463> A_IWL<6462> A_IWL<6461> A_IWL<6460> A_IWL<6459> A_IWL<6458> A_IWL<6457> A_IWL<6456> A_IWL<6455> A_IWL<6454> A_IWL<6453> A_IWL<6452> A_IWL<6451> A_IWL<6450> A_IWL<6449> A_IWL<6448> A_IWL<6447> A_IWL<6446> A_IWL<6445> A_IWL<6444> A_IWL<6443> A_IWL<6442> A_IWL<6441> A_IWL<6440> A_IWL<6439> A_IWL<6438> A_IWL<6437> A_IWL<6436> A_IWL<6435> A_IWL<6434> A_IWL<6433> A_IWL<6432> A_IWL<6431> A_IWL<6430> A_IWL<6429> A_IWL<6428> A_IWL<6427> A_IWL<6426> A_IWL<6425> A_IWL<6424> A_IWL<6423> A_IWL<6422> A_IWL<6421> A_IWL<6420> A_IWL<6419> A_IWL<6418> A_IWL<6417> A_IWL<6416> A_IWL<6415> A_IWL<6414> A_IWL<6413> A_IWL<6412> A_IWL<6411> A_IWL<6410> A_IWL<6409> A_IWL<6408> A_IWL<6407> A_IWL<6406> A_IWL<6405> A_IWL<6404> A_IWL<6403> A_IWL<6402> A_IWL<6401> A_IWL<6400> A_IWL<6911> A_IWL<6910> A_IWL<6909> A_IWL<6908> A_IWL<6907> A_IWL<6906> A_IWL<6905> A_IWL<6904> A_IWL<6903> A_IWL<6902> A_IWL<6901> A_IWL<6900> A_IWL<6899> A_IWL<6898> A_IWL<6897> A_IWL<6896> A_IWL<6895> A_IWL<6894> A_IWL<6893> A_IWL<6892> A_IWL<6891> A_IWL<6890> A_IWL<6889> A_IWL<6888> A_IWL<6887> A_IWL<6886> A_IWL<6885> A_IWL<6884> A_IWL<6883> A_IWL<6882> A_IWL<6881> A_IWL<6880> A_IWL<6879> A_IWL<6878> A_IWL<6877> A_IWL<6876> A_IWL<6875> A_IWL<6874> A_IWL<6873> A_IWL<6872> A_IWL<6871> A_IWL<6870> A_IWL<6869> A_IWL<6868> A_IWL<6867> A_IWL<6866> A_IWL<6865> A_IWL<6864> A_IWL<6863> A_IWL<6862> A_IWL<6861> A_IWL<6860> A_IWL<6859> A_IWL<6858> A_IWL<6857> A_IWL<6856> A_IWL<6855> A_IWL<6854> A_IWL<6853> A_IWL<6852> A_IWL<6851> A_IWL<6850> A_IWL<6849> A_IWL<6848> A_IWL<6847> A_IWL<6846> A_IWL<6845> A_IWL<6844> A_IWL<6843> A_IWL<6842> A_IWL<6841> A_IWL<6840> A_IWL<6839> A_IWL<6838> A_IWL<6837> A_IWL<6836> A_IWL<6835> A_IWL<6834> A_IWL<6833> A_IWL<6832> A_IWL<6831> A_IWL<6830> A_IWL<6829> A_IWL<6828> A_IWL<6827> A_IWL<6826> A_IWL<6825> A_IWL<6824> A_IWL<6823> A_IWL<6822> A_IWL<6821> A_IWL<6820> A_IWL<6819> A_IWL<6818> A_IWL<6817> A_IWL<6816> A_IWL<6815> A_IWL<6814> A_IWL<6813> A_IWL<6812> A_IWL<6811> A_IWL<6810> A_IWL<6809> A_IWL<6808> A_IWL<6807> A_IWL<6806> A_IWL<6805> A_IWL<6804> A_IWL<6803> A_IWL<6802> A_IWL<6801> A_IWL<6800> A_IWL<6799> A_IWL<6798> A_IWL<6797> A_IWL<6796> A_IWL<6795> A_IWL<6794> A_IWL<6793> A_IWL<6792> A_IWL<6791> A_IWL<6790> A_IWL<6789> A_IWL<6788> A_IWL<6787> A_IWL<6786> A_IWL<6785> A_IWL<6784> A_IWL<6783> A_IWL<6782> A_IWL<6781> A_IWL<6780> A_IWL<6779> A_IWL<6778> A_IWL<6777> A_IWL<6776> A_IWL<6775> A_IWL<6774> A_IWL<6773> A_IWL<6772> A_IWL<6771> A_IWL<6770> A_IWL<6769> A_IWL<6768> A_IWL<6767> A_IWL<6766> A_IWL<6765> A_IWL<6764> A_IWL<6763> A_IWL<6762> A_IWL<6761> A_IWL<6760> A_IWL<6759> A_IWL<6758> A_IWL<6757> A_IWL<6756> A_IWL<6755> A_IWL<6754> A_IWL<6753> A_IWL<6752> A_IWL<6751> A_IWL<6750> A_IWL<6749> A_IWL<6748> A_IWL<6747> A_IWL<6746> A_IWL<6745> A_IWL<6744> A_IWL<6743> A_IWL<6742> A_IWL<6741> A_IWL<6740> A_IWL<6739> A_IWL<6738> A_IWL<6737> A_IWL<6736> A_IWL<6735> A_IWL<6734> A_IWL<6733> A_IWL<6732> A_IWL<6731> A_IWL<6730> A_IWL<6729> A_IWL<6728> A_IWL<6727> A_IWL<6726> A_IWL<6725> A_IWL<6724> A_IWL<6723> A_IWL<6722> A_IWL<6721> A_IWL<6720> A_IWL<6719> A_IWL<6718> A_IWL<6717> A_IWL<6716> A_IWL<6715> A_IWL<6714> A_IWL<6713> A_IWL<6712> A_IWL<6711> A_IWL<6710> A_IWL<6709> A_IWL<6708> A_IWL<6707> A_IWL<6706> A_IWL<6705> A_IWL<6704> A_IWL<6703> A_IWL<6702> A_IWL<6701> A_IWL<6700> A_IWL<6699> A_IWL<6698> A_IWL<6697> A_IWL<6696> A_IWL<6695> A_IWL<6694> A_IWL<6693> A_IWL<6692> A_IWL<6691> A_IWL<6690> A_IWL<6689> A_IWL<6688> A_IWL<6687> A_IWL<6686> A_IWL<6685> A_IWL<6684> A_IWL<6683> A_IWL<6682> A_IWL<6681> A_IWL<6680> A_IWL<6679> A_IWL<6678> A_IWL<6677> A_IWL<6676> A_IWL<6675> A_IWL<6674> A_IWL<6673> A_IWL<6672> A_IWL<6671> A_IWL<6670> A_IWL<6669> A_IWL<6668> A_IWL<6667> A_IWL<6666> A_IWL<6665> A_IWL<6664> A_IWL<6663> A_IWL<6662> A_IWL<6661> A_IWL<6660> A_IWL<6659> A_IWL<6658> A_IWL<6657> A_IWL<6656> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<25> A_BLC<51> A_BLC<50> A_BLC_TOP<51> A_BLC_TOP<50> A_BLT<51> A_BLT<50> A_BLT_TOP<51> A_BLT_TOP<50> A_IWL<6399> A_IWL<6398> A_IWL<6397> A_IWL<6396> A_IWL<6395> A_IWL<6394> A_IWL<6393> A_IWL<6392> A_IWL<6391> A_IWL<6390> A_IWL<6389> A_IWL<6388> A_IWL<6387> A_IWL<6386> A_IWL<6385> A_IWL<6384> A_IWL<6383> A_IWL<6382> A_IWL<6381> A_IWL<6380> A_IWL<6379> A_IWL<6378> A_IWL<6377> A_IWL<6376> A_IWL<6375> A_IWL<6374> A_IWL<6373> A_IWL<6372> A_IWL<6371> A_IWL<6370> A_IWL<6369> A_IWL<6368> A_IWL<6367> A_IWL<6366> A_IWL<6365> A_IWL<6364> A_IWL<6363> A_IWL<6362> A_IWL<6361> A_IWL<6360> A_IWL<6359> A_IWL<6358> A_IWL<6357> A_IWL<6356> A_IWL<6355> A_IWL<6354> A_IWL<6353> A_IWL<6352> A_IWL<6351> A_IWL<6350> A_IWL<6349> A_IWL<6348> A_IWL<6347> A_IWL<6346> A_IWL<6345> A_IWL<6344> A_IWL<6343> A_IWL<6342> A_IWL<6341> A_IWL<6340> A_IWL<6339> A_IWL<6338> A_IWL<6337> A_IWL<6336> A_IWL<6335> A_IWL<6334> A_IWL<6333> A_IWL<6332> A_IWL<6331> A_IWL<6330> A_IWL<6329> A_IWL<6328> A_IWL<6327> A_IWL<6326> A_IWL<6325> A_IWL<6324> A_IWL<6323> A_IWL<6322> A_IWL<6321> A_IWL<6320> A_IWL<6319> A_IWL<6318> A_IWL<6317> A_IWL<6316> A_IWL<6315> A_IWL<6314> A_IWL<6313> A_IWL<6312> A_IWL<6311> A_IWL<6310> A_IWL<6309> A_IWL<6308> A_IWL<6307> A_IWL<6306> A_IWL<6305> A_IWL<6304> A_IWL<6303> A_IWL<6302> A_IWL<6301> A_IWL<6300> A_IWL<6299> A_IWL<6298> A_IWL<6297> A_IWL<6296> A_IWL<6295> A_IWL<6294> A_IWL<6293> A_IWL<6292> A_IWL<6291> A_IWL<6290> A_IWL<6289> A_IWL<6288> A_IWL<6287> A_IWL<6286> A_IWL<6285> A_IWL<6284> A_IWL<6283> A_IWL<6282> A_IWL<6281> A_IWL<6280> A_IWL<6279> A_IWL<6278> A_IWL<6277> A_IWL<6276> A_IWL<6275> A_IWL<6274> A_IWL<6273> A_IWL<6272> A_IWL<6271> A_IWL<6270> A_IWL<6269> A_IWL<6268> A_IWL<6267> A_IWL<6266> A_IWL<6265> A_IWL<6264> A_IWL<6263> A_IWL<6262> A_IWL<6261> A_IWL<6260> A_IWL<6259> A_IWL<6258> A_IWL<6257> A_IWL<6256> A_IWL<6255> A_IWL<6254> A_IWL<6253> A_IWL<6252> A_IWL<6251> A_IWL<6250> A_IWL<6249> A_IWL<6248> A_IWL<6247> A_IWL<6246> A_IWL<6245> A_IWL<6244> A_IWL<6243> A_IWL<6242> A_IWL<6241> A_IWL<6240> A_IWL<6239> A_IWL<6238> A_IWL<6237> A_IWL<6236> A_IWL<6235> A_IWL<6234> A_IWL<6233> A_IWL<6232> A_IWL<6231> A_IWL<6230> A_IWL<6229> A_IWL<6228> A_IWL<6227> A_IWL<6226> A_IWL<6225> A_IWL<6224> A_IWL<6223> A_IWL<6222> A_IWL<6221> A_IWL<6220> A_IWL<6219> A_IWL<6218> A_IWL<6217> A_IWL<6216> A_IWL<6215> A_IWL<6214> A_IWL<6213> A_IWL<6212> A_IWL<6211> A_IWL<6210> A_IWL<6209> A_IWL<6208> A_IWL<6207> A_IWL<6206> A_IWL<6205> A_IWL<6204> A_IWL<6203> A_IWL<6202> A_IWL<6201> A_IWL<6200> A_IWL<6199> A_IWL<6198> A_IWL<6197> A_IWL<6196> A_IWL<6195> A_IWL<6194> A_IWL<6193> A_IWL<6192> A_IWL<6191> A_IWL<6190> A_IWL<6189> A_IWL<6188> A_IWL<6187> A_IWL<6186> A_IWL<6185> A_IWL<6184> A_IWL<6183> A_IWL<6182> A_IWL<6181> A_IWL<6180> A_IWL<6179> A_IWL<6178> A_IWL<6177> A_IWL<6176> A_IWL<6175> A_IWL<6174> A_IWL<6173> A_IWL<6172> A_IWL<6171> A_IWL<6170> A_IWL<6169> A_IWL<6168> A_IWL<6167> A_IWL<6166> A_IWL<6165> A_IWL<6164> A_IWL<6163> A_IWL<6162> A_IWL<6161> A_IWL<6160> A_IWL<6159> A_IWL<6158> A_IWL<6157> A_IWL<6156> A_IWL<6155> A_IWL<6154> A_IWL<6153> A_IWL<6152> A_IWL<6151> A_IWL<6150> A_IWL<6149> A_IWL<6148> A_IWL<6147> A_IWL<6146> A_IWL<6145> A_IWL<6144> A_IWL<6655> A_IWL<6654> A_IWL<6653> A_IWL<6652> A_IWL<6651> A_IWL<6650> A_IWL<6649> A_IWL<6648> A_IWL<6647> A_IWL<6646> A_IWL<6645> A_IWL<6644> A_IWL<6643> A_IWL<6642> A_IWL<6641> A_IWL<6640> A_IWL<6639> A_IWL<6638> A_IWL<6637> A_IWL<6636> A_IWL<6635> A_IWL<6634> A_IWL<6633> A_IWL<6632> A_IWL<6631> A_IWL<6630> A_IWL<6629> A_IWL<6628> A_IWL<6627> A_IWL<6626> A_IWL<6625> A_IWL<6624> A_IWL<6623> A_IWL<6622> A_IWL<6621> A_IWL<6620> A_IWL<6619> A_IWL<6618> A_IWL<6617> A_IWL<6616> A_IWL<6615> A_IWL<6614> A_IWL<6613> A_IWL<6612> A_IWL<6611> A_IWL<6610> A_IWL<6609> A_IWL<6608> A_IWL<6607> A_IWL<6606> A_IWL<6605> A_IWL<6604> A_IWL<6603> A_IWL<6602> A_IWL<6601> A_IWL<6600> A_IWL<6599> A_IWL<6598> A_IWL<6597> A_IWL<6596> A_IWL<6595> A_IWL<6594> A_IWL<6593> A_IWL<6592> A_IWL<6591> A_IWL<6590> A_IWL<6589> A_IWL<6588> A_IWL<6587> A_IWL<6586> A_IWL<6585> A_IWL<6584> A_IWL<6583> A_IWL<6582> A_IWL<6581> A_IWL<6580> A_IWL<6579> A_IWL<6578> A_IWL<6577> A_IWL<6576> A_IWL<6575> A_IWL<6574> A_IWL<6573> A_IWL<6572> A_IWL<6571> A_IWL<6570> A_IWL<6569> A_IWL<6568> A_IWL<6567> A_IWL<6566> A_IWL<6565> A_IWL<6564> A_IWL<6563> A_IWL<6562> A_IWL<6561> A_IWL<6560> A_IWL<6559> A_IWL<6558> A_IWL<6557> A_IWL<6556> A_IWL<6555> A_IWL<6554> A_IWL<6553> A_IWL<6552> A_IWL<6551> A_IWL<6550> A_IWL<6549> A_IWL<6548> A_IWL<6547> A_IWL<6546> A_IWL<6545> A_IWL<6544> A_IWL<6543> A_IWL<6542> A_IWL<6541> A_IWL<6540> A_IWL<6539> A_IWL<6538> A_IWL<6537> A_IWL<6536> A_IWL<6535> A_IWL<6534> A_IWL<6533> A_IWL<6532> A_IWL<6531> A_IWL<6530> A_IWL<6529> A_IWL<6528> A_IWL<6527> A_IWL<6526> A_IWL<6525> A_IWL<6524> A_IWL<6523> A_IWL<6522> A_IWL<6521> A_IWL<6520> A_IWL<6519> A_IWL<6518> A_IWL<6517> A_IWL<6516> A_IWL<6515> A_IWL<6514> A_IWL<6513> A_IWL<6512> A_IWL<6511> A_IWL<6510> A_IWL<6509> A_IWL<6508> A_IWL<6507> A_IWL<6506> A_IWL<6505> A_IWL<6504> A_IWL<6503> A_IWL<6502> A_IWL<6501> A_IWL<6500> A_IWL<6499> A_IWL<6498> A_IWL<6497> A_IWL<6496> A_IWL<6495> A_IWL<6494> A_IWL<6493> A_IWL<6492> A_IWL<6491> A_IWL<6490> A_IWL<6489> A_IWL<6488> A_IWL<6487> A_IWL<6486> A_IWL<6485> A_IWL<6484> A_IWL<6483> A_IWL<6482> A_IWL<6481> A_IWL<6480> A_IWL<6479> A_IWL<6478> A_IWL<6477> A_IWL<6476> A_IWL<6475> A_IWL<6474> A_IWL<6473> A_IWL<6472> A_IWL<6471> A_IWL<6470> A_IWL<6469> A_IWL<6468> A_IWL<6467> A_IWL<6466> A_IWL<6465> A_IWL<6464> A_IWL<6463> A_IWL<6462> A_IWL<6461> A_IWL<6460> A_IWL<6459> A_IWL<6458> A_IWL<6457> A_IWL<6456> A_IWL<6455> A_IWL<6454> A_IWL<6453> A_IWL<6452> A_IWL<6451> A_IWL<6450> A_IWL<6449> A_IWL<6448> A_IWL<6447> A_IWL<6446> A_IWL<6445> A_IWL<6444> A_IWL<6443> A_IWL<6442> A_IWL<6441> A_IWL<6440> A_IWL<6439> A_IWL<6438> A_IWL<6437> A_IWL<6436> A_IWL<6435> A_IWL<6434> A_IWL<6433> A_IWL<6432> A_IWL<6431> A_IWL<6430> A_IWL<6429> A_IWL<6428> A_IWL<6427> A_IWL<6426> A_IWL<6425> A_IWL<6424> A_IWL<6423> A_IWL<6422> A_IWL<6421> A_IWL<6420> A_IWL<6419> A_IWL<6418> A_IWL<6417> A_IWL<6416> A_IWL<6415> A_IWL<6414> A_IWL<6413> A_IWL<6412> A_IWL<6411> A_IWL<6410> A_IWL<6409> A_IWL<6408> A_IWL<6407> A_IWL<6406> A_IWL<6405> A_IWL<6404> A_IWL<6403> A_IWL<6402> A_IWL<6401> A_IWL<6400> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<24> A_BLC<49> A_BLC<48> A_BLC_TOP<49> A_BLC_TOP<48> A_BLT<49> A_BLT<48> A_BLT_TOP<49> A_BLT_TOP<48> A_IWL<6143> A_IWL<6142> A_IWL<6141> A_IWL<6140> A_IWL<6139> A_IWL<6138> A_IWL<6137> A_IWL<6136> A_IWL<6135> A_IWL<6134> A_IWL<6133> A_IWL<6132> A_IWL<6131> A_IWL<6130> A_IWL<6129> A_IWL<6128> A_IWL<6127> A_IWL<6126> A_IWL<6125> A_IWL<6124> A_IWL<6123> A_IWL<6122> A_IWL<6121> A_IWL<6120> A_IWL<6119> A_IWL<6118> A_IWL<6117> A_IWL<6116> A_IWL<6115> A_IWL<6114> A_IWL<6113> A_IWL<6112> A_IWL<6111> A_IWL<6110> A_IWL<6109> A_IWL<6108> A_IWL<6107> A_IWL<6106> A_IWL<6105> A_IWL<6104> A_IWL<6103> A_IWL<6102> A_IWL<6101> A_IWL<6100> A_IWL<6099> A_IWL<6098> A_IWL<6097> A_IWL<6096> A_IWL<6095> A_IWL<6094> A_IWL<6093> A_IWL<6092> A_IWL<6091> A_IWL<6090> A_IWL<6089> A_IWL<6088> A_IWL<6087> A_IWL<6086> A_IWL<6085> A_IWL<6084> A_IWL<6083> A_IWL<6082> A_IWL<6081> A_IWL<6080> A_IWL<6079> A_IWL<6078> A_IWL<6077> A_IWL<6076> A_IWL<6075> A_IWL<6074> A_IWL<6073> A_IWL<6072> A_IWL<6071> A_IWL<6070> A_IWL<6069> A_IWL<6068> A_IWL<6067> A_IWL<6066> A_IWL<6065> A_IWL<6064> A_IWL<6063> A_IWL<6062> A_IWL<6061> A_IWL<6060> A_IWL<6059> A_IWL<6058> A_IWL<6057> A_IWL<6056> A_IWL<6055> A_IWL<6054> A_IWL<6053> A_IWL<6052> A_IWL<6051> A_IWL<6050> A_IWL<6049> A_IWL<6048> A_IWL<6047> A_IWL<6046> A_IWL<6045> A_IWL<6044> A_IWL<6043> A_IWL<6042> A_IWL<6041> A_IWL<6040> A_IWL<6039> A_IWL<6038> A_IWL<6037> A_IWL<6036> A_IWL<6035> A_IWL<6034> A_IWL<6033> A_IWL<6032> A_IWL<6031> A_IWL<6030> A_IWL<6029> A_IWL<6028> A_IWL<6027> A_IWL<6026> A_IWL<6025> A_IWL<6024> A_IWL<6023> A_IWL<6022> A_IWL<6021> A_IWL<6020> A_IWL<6019> A_IWL<6018> A_IWL<6017> A_IWL<6016> A_IWL<6015> A_IWL<6014> A_IWL<6013> A_IWL<6012> A_IWL<6011> A_IWL<6010> A_IWL<6009> A_IWL<6008> A_IWL<6007> A_IWL<6006> A_IWL<6005> A_IWL<6004> A_IWL<6003> A_IWL<6002> A_IWL<6001> A_IWL<6000> A_IWL<5999> A_IWL<5998> A_IWL<5997> A_IWL<5996> A_IWL<5995> A_IWL<5994> A_IWL<5993> A_IWL<5992> A_IWL<5991> A_IWL<5990> A_IWL<5989> A_IWL<5988> A_IWL<5987> A_IWL<5986> A_IWL<5985> A_IWL<5984> A_IWL<5983> A_IWL<5982> A_IWL<5981> A_IWL<5980> A_IWL<5979> A_IWL<5978> A_IWL<5977> A_IWL<5976> A_IWL<5975> A_IWL<5974> A_IWL<5973> A_IWL<5972> A_IWL<5971> A_IWL<5970> A_IWL<5969> A_IWL<5968> A_IWL<5967> A_IWL<5966> A_IWL<5965> A_IWL<5964> A_IWL<5963> A_IWL<5962> A_IWL<5961> A_IWL<5960> A_IWL<5959> A_IWL<5958> A_IWL<5957> A_IWL<5956> A_IWL<5955> A_IWL<5954> A_IWL<5953> A_IWL<5952> A_IWL<5951> A_IWL<5950> A_IWL<5949> A_IWL<5948> A_IWL<5947> A_IWL<5946> A_IWL<5945> A_IWL<5944> A_IWL<5943> A_IWL<5942> A_IWL<5941> A_IWL<5940> A_IWL<5939> A_IWL<5938> A_IWL<5937> A_IWL<5936> A_IWL<5935> A_IWL<5934> A_IWL<5933> A_IWL<5932> A_IWL<5931> A_IWL<5930> A_IWL<5929> A_IWL<5928> A_IWL<5927> A_IWL<5926> A_IWL<5925> A_IWL<5924> A_IWL<5923> A_IWL<5922> A_IWL<5921> A_IWL<5920> A_IWL<5919> A_IWL<5918> A_IWL<5917> A_IWL<5916> A_IWL<5915> A_IWL<5914> A_IWL<5913> A_IWL<5912> A_IWL<5911> A_IWL<5910> A_IWL<5909> A_IWL<5908> A_IWL<5907> A_IWL<5906> A_IWL<5905> A_IWL<5904> A_IWL<5903> A_IWL<5902> A_IWL<5901> A_IWL<5900> A_IWL<5899> A_IWL<5898> A_IWL<5897> A_IWL<5896> A_IWL<5895> A_IWL<5894> A_IWL<5893> A_IWL<5892> A_IWL<5891> A_IWL<5890> A_IWL<5889> A_IWL<5888> A_IWL<6399> A_IWL<6398> A_IWL<6397> A_IWL<6396> A_IWL<6395> A_IWL<6394> A_IWL<6393> A_IWL<6392> A_IWL<6391> A_IWL<6390> A_IWL<6389> A_IWL<6388> A_IWL<6387> A_IWL<6386> A_IWL<6385> A_IWL<6384> A_IWL<6383> A_IWL<6382> A_IWL<6381> A_IWL<6380> A_IWL<6379> A_IWL<6378> A_IWL<6377> A_IWL<6376> A_IWL<6375> A_IWL<6374> A_IWL<6373> A_IWL<6372> A_IWL<6371> A_IWL<6370> A_IWL<6369> A_IWL<6368> A_IWL<6367> A_IWL<6366> A_IWL<6365> A_IWL<6364> A_IWL<6363> A_IWL<6362> A_IWL<6361> A_IWL<6360> A_IWL<6359> A_IWL<6358> A_IWL<6357> A_IWL<6356> A_IWL<6355> A_IWL<6354> A_IWL<6353> A_IWL<6352> A_IWL<6351> A_IWL<6350> A_IWL<6349> A_IWL<6348> A_IWL<6347> A_IWL<6346> A_IWL<6345> A_IWL<6344> A_IWL<6343> A_IWL<6342> A_IWL<6341> A_IWL<6340> A_IWL<6339> A_IWL<6338> A_IWL<6337> A_IWL<6336> A_IWL<6335> A_IWL<6334> A_IWL<6333> A_IWL<6332> A_IWL<6331> A_IWL<6330> A_IWL<6329> A_IWL<6328> A_IWL<6327> A_IWL<6326> A_IWL<6325> A_IWL<6324> A_IWL<6323> A_IWL<6322> A_IWL<6321> A_IWL<6320> A_IWL<6319> A_IWL<6318> A_IWL<6317> A_IWL<6316> A_IWL<6315> A_IWL<6314> A_IWL<6313> A_IWL<6312> A_IWL<6311> A_IWL<6310> A_IWL<6309> A_IWL<6308> A_IWL<6307> A_IWL<6306> A_IWL<6305> A_IWL<6304> A_IWL<6303> A_IWL<6302> A_IWL<6301> A_IWL<6300> A_IWL<6299> A_IWL<6298> A_IWL<6297> A_IWL<6296> A_IWL<6295> A_IWL<6294> A_IWL<6293> A_IWL<6292> A_IWL<6291> A_IWL<6290> A_IWL<6289> A_IWL<6288> A_IWL<6287> A_IWL<6286> A_IWL<6285> A_IWL<6284> A_IWL<6283> A_IWL<6282> A_IWL<6281> A_IWL<6280> A_IWL<6279> A_IWL<6278> A_IWL<6277> A_IWL<6276> A_IWL<6275> A_IWL<6274> A_IWL<6273> A_IWL<6272> A_IWL<6271> A_IWL<6270> A_IWL<6269> A_IWL<6268> A_IWL<6267> A_IWL<6266> A_IWL<6265> A_IWL<6264> A_IWL<6263> A_IWL<6262> A_IWL<6261> A_IWL<6260> A_IWL<6259> A_IWL<6258> A_IWL<6257> A_IWL<6256> A_IWL<6255> A_IWL<6254> A_IWL<6253> A_IWL<6252> A_IWL<6251> A_IWL<6250> A_IWL<6249> A_IWL<6248> A_IWL<6247> A_IWL<6246> A_IWL<6245> A_IWL<6244> A_IWL<6243> A_IWL<6242> A_IWL<6241> A_IWL<6240> A_IWL<6239> A_IWL<6238> A_IWL<6237> A_IWL<6236> A_IWL<6235> A_IWL<6234> A_IWL<6233> A_IWL<6232> A_IWL<6231> A_IWL<6230> A_IWL<6229> A_IWL<6228> A_IWL<6227> A_IWL<6226> A_IWL<6225> A_IWL<6224> A_IWL<6223> A_IWL<6222> A_IWL<6221> A_IWL<6220> A_IWL<6219> A_IWL<6218> A_IWL<6217> A_IWL<6216> A_IWL<6215> A_IWL<6214> A_IWL<6213> A_IWL<6212> A_IWL<6211> A_IWL<6210> A_IWL<6209> A_IWL<6208> A_IWL<6207> A_IWL<6206> A_IWL<6205> A_IWL<6204> A_IWL<6203> A_IWL<6202> A_IWL<6201> A_IWL<6200> A_IWL<6199> A_IWL<6198> A_IWL<6197> A_IWL<6196> A_IWL<6195> A_IWL<6194> A_IWL<6193> A_IWL<6192> A_IWL<6191> A_IWL<6190> A_IWL<6189> A_IWL<6188> A_IWL<6187> A_IWL<6186> A_IWL<6185> A_IWL<6184> A_IWL<6183> A_IWL<6182> A_IWL<6181> A_IWL<6180> A_IWL<6179> A_IWL<6178> A_IWL<6177> A_IWL<6176> A_IWL<6175> A_IWL<6174> A_IWL<6173> A_IWL<6172> A_IWL<6171> A_IWL<6170> A_IWL<6169> A_IWL<6168> A_IWL<6167> A_IWL<6166> A_IWL<6165> A_IWL<6164> A_IWL<6163> A_IWL<6162> A_IWL<6161> A_IWL<6160> A_IWL<6159> A_IWL<6158> A_IWL<6157> A_IWL<6156> A_IWL<6155> A_IWL<6154> A_IWL<6153> A_IWL<6152> A_IWL<6151> A_IWL<6150> A_IWL<6149> A_IWL<6148> A_IWL<6147> A_IWL<6146> A_IWL<6145> A_IWL<6144> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<23> A_BLC<47> A_BLC<46> A_BLC_TOP<47> A_BLC_TOP<46> A_BLT<47> A_BLT<46> A_BLT_TOP<47> A_BLT_TOP<46> A_IWL<5887> A_IWL<5886> A_IWL<5885> A_IWL<5884> A_IWL<5883> A_IWL<5882> A_IWL<5881> A_IWL<5880> A_IWL<5879> A_IWL<5878> A_IWL<5877> A_IWL<5876> A_IWL<5875> A_IWL<5874> A_IWL<5873> A_IWL<5872> A_IWL<5871> A_IWL<5870> A_IWL<5869> A_IWL<5868> A_IWL<5867> A_IWL<5866> A_IWL<5865> A_IWL<5864> A_IWL<5863> A_IWL<5862> A_IWL<5861> A_IWL<5860> A_IWL<5859> A_IWL<5858> A_IWL<5857> A_IWL<5856> A_IWL<5855> A_IWL<5854> A_IWL<5853> A_IWL<5852> A_IWL<5851> A_IWL<5850> A_IWL<5849> A_IWL<5848> A_IWL<5847> A_IWL<5846> A_IWL<5845> A_IWL<5844> A_IWL<5843> A_IWL<5842> A_IWL<5841> A_IWL<5840> A_IWL<5839> A_IWL<5838> A_IWL<5837> A_IWL<5836> A_IWL<5835> A_IWL<5834> A_IWL<5833> A_IWL<5832> A_IWL<5831> A_IWL<5830> A_IWL<5829> A_IWL<5828> A_IWL<5827> A_IWL<5826> A_IWL<5825> A_IWL<5824> A_IWL<5823> A_IWL<5822> A_IWL<5821> A_IWL<5820> A_IWL<5819> A_IWL<5818> A_IWL<5817> A_IWL<5816> A_IWL<5815> A_IWL<5814> A_IWL<5813> A_IWL<5812> A_IWL<5811> A_IWL<5810> A_IWL<5809> A_IWL<5808> A_IWL<5807> A_IWL<5806> A_IWL<5805> A_IWL<5804> A_IWL<5803> A_IWL<5802> A_IWL<5801> A_IWL<5800> A_IWL<5799> A_IWL<5798> A_IWL<5797> A_IWL<5796> A_IWL<5795> A_IWL<5794> A_IWL<5793> A_IWL<5792> A_IWL<5791> A_IWL<5790> A_IWL<5789> A_IWL<5788> A_IWL<5787> A_IWL<5786> A_IWL<5785> A_IWL<5784> A_IWL<5783> A_IWL<5782> A_IWL<5781> A_IWL<5780> A_IWL<5779> A_IWL<5778> A_IWL<5777> A_IWL<5776> A_IWL<5775> A_IWL<5774> A_IWL<5773> A_IWL<5772> A_IWL<5771> A_IWL<5770> A_IWL<5769> A_IWL<5768> A_IWL<5767> A_IWL<5766> A_IWL<5765> A_IWL<5764> A_IWL<5763> A_IWL<5762> A_IWL<5761> A_IWL<5760> A_IWL<5759> A_IWL<5758> A_IWL<5757> A_IWL<5756> A_IWL<5755> A_IWL<5754> A_IWL<5753> A_IWL<5752> A_IWL<5751> A_IWL<5750> A_IWL<5749> A_IWL<5748> A_IWL<5747> A_IWL<5746> A_IWL<5745> A_IWL<5744> A_IWL<5743> A_IWL<5742> A_IWL<5741> A_IWL<5740> A_IWL<5739> A_IWL<5738> A_IWL<5737> A_IWL<5736> A_IWL<5735> A_IWL<5734> A_IWL<5733> A_IWL<5732> A_IWL<5731> A_IWL<5730> A_IWL<5729> A_IWL<5728> A_IWL<5727> A_IWL<5726> A_IWL<5725> A_IWL<5724> A_IWL<5723> A_IWL<5722> A_IWL<5721> A_IWL<5720> A_IWL<5719> A_IWL<5718> A_IWL<5717> A_IWL<5716> A_IWL<5715> A_IWL<5714> A_IWL<5713> A_IWL<5712> A_IWL<5711> A_IWL<5710> A_IWL<5709> A_IWL<5708> A_IWL<5707> A_IWL<5706> A_IWL<5705> A_IWL<5704> A_IWL<5703> A_IWL<5702> A_IWL<5701> A_IWL<5700> A_IWL<5699> A_IWL<5698> A_IWL<5697> A_IWL<5696> A_IWL<5695> A_IWL<5694> A_IWL<5693> A_IWL<5692> A_IWL<5691> A_IWL<5690> A_IWL<5689> A_IWL<5688> A_IWL<5687> A_IWL<5686> A_IWL<5685> A_IWL<5684> A_IWL<5683> A_IWL<5682> A_IWL<5681> A_IWL<5680> A_IWL<5679> A_IWL<5678> A_IWL<5677> A_IWL<5676> A_IWL<5675> A_IWL<5674> A_IWL<5673> A_IWL<5672> A_IWL<5671> A_IWL<5670> A_IWL<5669> A_IWL<5668> A_IWL<5667> A_IWL<5666> A_IWL<5665> A_IWL<5664> A_IWL<5663> A_IWL<5662> A_IWL<5661> A_IWL<5660> A_IWL<5659> A_IWL<5658> A_IWL<5657> A_IWL<5656> A_IWL<5655> A_IWL<5654> A_IWL<5653> A_IWL<5652> A_IWL<5651> A_IWL<5650> A_IWL<5649> A_IWL<5648> A_IWL<5647> A_IWL<5646> A_IWL<5645> A_IWL<5644> A_IWL<5643> A_IWL<5642> A_IWL<5641> A_IWL<5640> A_IWL<5639> A_IWL<5638> A_IWL<5637> A_IWL<5636> A_IWL<5635> A_IWL<5634> A_IWL<5633> A_IWL<5632> A_IWL<6143> A_IWL<6142> A_IWL<6141> A_IWL<6140> A_IWL<6139> A_IWL<6138> A_IWL<6137> A_IWL<6136> A_IWL<6135> A_IWL<6134> A_IWL<6133> A_IWL<6132> A_IWL<6131> A_IWL<6130> A_IWL<6129> A_IWL<6128> A_IWL<6127> A_IWL<6126> A_IWL<6125> A_IWL<6124> A_IWL<6123> A_IWL<6122> A_IWL<6121> A_IWL<6120> A_IWL<6119> A_IWL<6118> A_IWL<6117> A_IWL<6116> A_IWL<6115> A_IWL<6114> A_IWL<6113> A_IWL<6112> A_IWL<6111> A_IWL<6110> A_IWL<6109> A_IWL<6108> A_IWL<6107> A_IWL<6106> A_IWL<6105> A_IWL<6104> A_IWL<6103> A_IWL<6102> A_IWL<6101> A_IWL<6100> A_IWL<6099> A_IWL<6098> A_IWL<6097> A_IWL<6096> A_IWL<6095> A_IWL<6094> A_IWL<6093> A_IWL<6092> A_IWL<6091> A_IWL<6090> A_IWL<6089> A_IWL<6088> A_IWL<6087> A_IWL<6086> A_IWL<6085> A_IWL<6084> A_IWL<6083> A_IWL<6082> A_IWL<6081> A_IWL<6080> A_IWL<6079> A_IWL<6078> A_IWL<6077> A_IWL<6076> A_IWL<6075> A_IWL<6074> A_IWL<6073> A_IWL<6072> A_IWL<6071> A_IWL<6070> A_IWL<6069> A_IWL<6068> A_IWL<6067> A_IWL<6066> A_IWL<6065> A_IWL<6064> A_IWL<6063> A_IWL<6062> A_IWL<6061> A_IWL<6060> A_IWL<6059> A_IWL<6058> A_IWL<6057> A_IWL<6056> A_IWL<6055> A_IWL<6054> A_IWL<6053> A_IWL<6052> A_IWL<6051> A_IWL<6050> A_IWL<6049> A_IWL<6048> A_IWL<6047> A_IWL<6046> A_IWL<6045> A_IWL<6044> A_IWL<6043> A_IWL<6042> A_IWL<6041> A_IWL<6040> A_IWL<6039> A_IWL<6038> A_IWL<6037> A_IWL<6036> A_IWL<6035> A_IWL<6034> A_IWL<6033> A_IWL<6032> A_IWL<6031> A_IWL<6030> A_IWL<6029> A_IWL<6028> A_IWL<6027> A_IWL<6026> A_IWL<6025> A_IWL<6024> A_IWL<6023> A_IWL<6022> A_IWL<6021> A_IWL<6020> A_IWL<6019> A_IWL<6018> A_IWL<6017> A_IWL<6016> A_IWL<6015> A_IWL<6014> A_IWL<6013> A_IWL<6012> A_IWL<6011> A_IWL<6010> A_IWL<6009> A_IWL<6008> A_IWL<6007> A_IWL<6006> A_IWL<6005> A_IWL<6004> A_IWL<6003> A_IWL<6002> A_IWL<6001> A_IWL<6000> A_IWL<5999> A_IWL<5998> A_IWL<5997> A_IWL<5996> A_IWL<5995> A_IWL<5994> A_IWL<5993> A_IWL<5992> A_IWL<5991> A_IWL<5990> A_IWL<5989> A_IWL<5988> A_IWL<5987> A_IWL<5986> A_IWL<5985> A_IWL<5984> A_IWL<5983> A_IWL<5982> A_IWL<5981> A_IWL<5980> A_IWL<5979> A_IWL<5978> A_IWL<5977> A_IWL<5976> A_IWL<5975> A_IWL<5974> A_IWL<5973> A_IWL<5972> A_IWL<5971> A_IWL<5970> A_IWL<5969> A_IWL<5968> A_IWL<5967> A_IWL<5966> A_IWL<5965> A_IWL<5964> A_IWL<5963> A_IWL<5962> A_IWL<5961> A_IWL<5960> A_IWL<5959> A_IWL<5958> A_IWL<5957> A_IWL<5956> A_IWL<5955> A_IWL<5954> A_IWL<5953> A_IWL<5952> A_IWL<5951> A_IWL<5950> A_IWL<5949> A_IWL<5948> A_IWL<5947> A_IWL<5946> A_IWL<5945> A_IWL<5944> A_IWL<5943> A_IWL<5942> A_IWL<5941> A_IWL<5940> A_IWL<5939> A_IWL<5938> A_IWL<5937> A_IWL<5936> A_IWL<5935> A_IWL<5934> A_IWL<5933> A_IWL<5932> A_IWL<5931> A_IWL<5930> A_IWL<5929> A_IWL<5928> A_IWL<5927> A_IWL<5926> A_IWL<5925> A_IWL<5924> A_IWL<5923> A_IWL<5922> A_IWL<5921> A_IWL<5920> A_IWL<5919> A_IWL<5918> A_IWL<5917> A_IWL<5916> A_IWL<5915> A_IWL<5914> A_IWL<5913> A_IWL<5912> A_IWL<5911> A_IWL<5910> A_IWL<5909> A_IWL<5908> A_IWL<5907> A_IWL<5906> A_IWL<5905> A_IWL<5904> A_IWL<5903> A_IWL<5902> A_IWL<5901> A_IWL<5900> A_IWL<5899> A_IWL<5898> A_IWL<5897> A_IWL<5896> A_IWL<5895> A_IWL<5894> A_IWL<5893> A_IWL<5892> A_IWL<5891> A_IWL<5890> A_IWL<5889> A_IWL<5888> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<22> A_BLC<45> A_BLC<44> A_BLC_TOP<45> A_BLC_TOP<44> A_BLT<45> A_BLT<44> A_BLT_TOP<45> A_BLT_TOP<44> A_IWL<5631> A_IWL<5630> A_IWL<5629> A_IWL<5628> A_IWL<5627> A_IWL<5626> A_IWL<5625> A_IWL<5624> A_IWL<5623> A_IWL<5622> A_IWL<5621> A_IWL<5620> A_IWL<5619> A_IWL<5618> A_IWL<5617> A_IWL<5616> A_IWL<5615> A_IWL<5614> A_IWL<5613> A_IWL<5612> A_IWL<5611> A_IWL<5610> A_IWL<5609> A_IWL<5608> A_IWL<5607> A_IWL<5606> A_IWL<5605> A_IWL<5604> A_IWL<5603> A_IWL<5602> A_IWL<5601> A_IWL<5600> A_IWL<5599> A_IWL<5598> A_IWL<5597> A_IWL<5596> A_IWL<5595> A_IWL<5594> A_IWL<5593> A_IWL<5592> A_IWL<5591> A_IWL<5590> A_IWL<5589> A_IWL<5588> A_IWL<5587> A_IWL<5586> A_IWL<5585> A_IWL<5584> A_IWL<5583> A_IWL<5582> A_IWL<5581> A_IWL<5580> A_IWL<5579> A_IWL<5578> A_IWL<5577> A_IWL<5576> A_IWL<5575> A_IWL<5574> A_IWL<5573> A_IWL<5572> A_IWL<5571> A_IWL<5570> A_IWL<5569> A_IWL<5568> A_IWL<5567> A_IWL<5566> A_IWL<5565> A_IWL<5564> A_IWL<5563> A_IWL<5562> A_IWL<5561> A_IWL<5560> A_IWL<5559> A_IWL<5558> A_IWL<5557> A_IWL<5556> A_IWL<5555> A_IWL<5554> A_IWL<5553> A_IWL<5552> A_IWL<5551> A_IWL<5550> A_IWL<5549> A_IWL<5548> A_IWL<5547> A_IWL<5546> A_IWL<5545> A_IWL<5544> A_IWL<5543> A_IWL<5542> A_IWL<5541> A_IWL<5540> A_IWL<5539> A_IWL<5538> A_IWL<5537> A_IWL<5536> A_IWL<5535> A_IWL<5534> A_IWL<5533> A_IWL<5532> A_IWL<5531> A_IWL<5530> A_IWL<5529> A_IWL<5528> A_IWL<5527> A_IWL<5526> A_IWL<5525> A_IWL<5524> A_IWL<5523> A_IWL<5522> A_IWL<5521> A_IWL<5520> A_IWL<5519> A_IWL<5518> A_IWL<5517> A_IWL<5516> A_IWL<5515> A_IWL<5514> A_IWL<5513> A_IWL<5512> A_IWL<5511> A_IWL<5510> A_IWL<5509> A_IWL<5508> A_IWL<5507> A_IWL<5506> A_IWL<5505> A_IWL<5504> A_IWL<5503> A_IWL<5502> A_IWL<5501> A_IWL<5500> A_IWL<5499> A_IWL<5498> A_IWL<5497> A_IWL<5496> A_IWL<5495> A_IWL<5494> A_IWL<5493> A_IWL<5492> A_IWL<5491> A_IWL<5490> A_IWL<5489> A_IWL<5488> A_IWL<5487> A_IWL<5486> A_IWL<5485> A_IWL<5484> A_IWL<5483> A_IWL<5482> A_IWL<5481> A_IWL<5480> A_IWL<5479> A_IWL<5478> A_IWL<5477> A_IWL<5476> A_IWL<5475> A_IWL<5474> A_IWL<5473> A_IWL<5472> A_IWL<5471> A_IWL<5470> A_IWL<5469> A_IWL<5468> A_IWL<5467> A_IWL<5466> A_IWL<5465> A_IWL<5464> A_IWL<5463> A_IWL<5462> A_IWL<5461> A_IWL<5460> A_IWL<5459> A_IWL<5458> A_IWL<5457> A_IWL<5456> A_IWL<5455> A_IWL<5454> A_IWL<5453> A_IWL<5452> A_IWL<5451> A_IWL<5450> A_IWL<5449> A_IWL<5448> A_IWL<5447> A_IWL<5446> A_IWL<5445> A_IWL<5444> A_IWL<5443> A_IWL<5442> A_IWL<5441> A_IWL<5440> A_IWL<5439> A_IWL<5438> A_IWL<5437> A_IWL<5436> A_IWL<5435> A_IWL<5434> A_IWL<5433> A_IWL<5432> A_IWL<5431> A_IWL<5430> A_IWL<5429> A_IWL<5428> A_IWL<5427> A_IWL<5426> A_IWL<5425> A_IWL<5424> A_IWL<5423> A_IWL<5422> A_IWL<5421> A_IWL<5420> A_IWL<5419> A_IWL<5418> A_IWL<5417> A_IWL<5416> A_IWL<5415> A_IWL<5414> A_IWL<5413> A_IWL<5412> A_IWL<5411> A_IWL<5410> A_IWL<5409> A_IWL<5408> A_IWL<5407> A_IWL<5406> A_IWL<5405> A_IWL<5404> A_IWL<5403> A_IWL<5402> A_IWL<5401> A_IWL<5400> A_IWL<5399> A_IWL<5398> A_IWL<5397> A_IWL<5396> A_IWL<5395> A_IWL<5394> A_IWL<5393> A_IWL<5392> A_IWL<5391> A_IWL<5390> A_IWL<5389> A_IWL<5388> A_IWL<5387> A_IWL<5386> A_IWL<5385> A_IWL<5384> A_IWL<5383> A_IWL<5382> A_IWL<5381> A_IWL<5380> A_IWL<5379> A_IWL<5378> A_IWL<5377> A_IWL<5376> A_IWL<5887> A_IWL<5886> A_IWL<5885> A_IWL<5884> A_IWL<5883> A_IWL<5882> A_IWL<5881> A_IWL<5880> A_IWL<5879> A_IWL<5878> A_IWL<5877> A_IWL<5876> A_IWL<5875> A_IWL<5874> A_IWL<5873> A_IWL<5872> A_IWL<5871> A_IWL<5870> A_IWL<5869> A_IWL<5868> A_IWL<5867> A_IWL<5866> A_IWL<5865> A_IWL<5864> A_IWL<5863> A_IWL<5862> A_IWL<5861> A_IWL<5860> A_IWL<5859> A_IWL<5858> A_IWL<5857> A_IWL<5856> A_IWL<5855> A_IWL<5854> A_IWL<5853> A_IWL<5852> A_IWL<5851> A_IWL<5850> A_IWL<5849> A_IWL<5848> A_IWL<5847> A_IWL<5846> A_IWL<5845> A_IWL<5844> A_IWL<5843> A_IWL<5842> A_IWL<5841> A_IWL<5840> A_IWL<5839> A_IWL<5838> A_IWL<5837> A_IWL<5836> A_IWL<5835> A_IWL<5834> A_IWL<5833> A_IWL<5832> A_IWL<5831> A_IWL<5830> A_IWL<5829> A_IWL<5828> A_IWL<5827> A_IWL<5826> A_IWL<5825> A_IWL<5824> A_IWL<5823> A_IWL<5822> A_IWL<5821> A_IWL<5820> A_IWL<5819> A_IWL<5818> A_IWL<5817> A_IWL<5816> A_IWL<5815> A_IWL<5814> A_IWL<5813> A_IWL<5812> A_IWL<5811> A_IWL<5810> A_IWL<5809> A_IWL<5808> A_IWL<5807> A_IWL<5806> A_IWL<5805> A_IWL<5804> A_IWL<5803> A_IWL<5802> A_IWL<5801> A_IWL<5800> A_IWL<5799> A_IWL<5798> A_IWL<5797> A_IWL<5796> A_IWL<5795> A_IWL<5794> A_IWL<5793> A_IWL<5792> A_IWL<5791> A_IWL<5790> A_IWL<5789> A_IWL<5788> A_IWL<5787> A_IWL<5786> A_IWL<5785> A_IWL<5784> A_IWL<5783> A_IWL<5782> A_IWL<5781> A_IWL<5780> A_IWL<5779> A_IWL<5778> A_IWL<5777> A_IWL<5776> A_IWL<5775> A_IWL<5774> A_IWL<5773> A_IWL<5772> A_IWL<5771> A_IWL<5770> A_IWL<5769> A_IWL<5768> A_IWL<5767> A_IWL<5766> A_IWL<5765> A_IWL<5764> A_IWL<5763> A_IWL<5762> A_IWL<5761> A_IWL<5760> A_IWL<5759> A_IWL<5758> A_IWL<5757> A_IWL<5756> A_IWL<5755> A_IWL<5754> A_IWL<5753> A_IWL<5752> A_IWL<5751> A_IWL<5750> A_IWL<5749> A_IWL<5748> A_IWL<5747> A_IWL<5746> A_IWL<5745> A_IWL<5744> A_IWL<5743> A_IWL<5742> A_IWL<5741> A_IWL<5740> A_IWL<5739> A_IWL<5738> A_IWL<5737> A_IWL<5736> A_IWL<5735> A_IWL<5734> A_IWL<5733> A_IWL<5732> A_IWL<5731> A_IWL<5730> A_IWL<5729> A_IWL<5728> A_IWL<5727> A_IWL<5726> A_IWL<5725> A_IWL<5724> A_IWL<5723> A_IWL<5722> A_IWL<5721> A_IWL<5720> A_IWL<5719> A_IWL<5718> A_IWL<5717> A_IWL<5716> A_IWL<5715> A_IWL<5714> A_IWL<5713> A_IWL<5712> A_IWL<5711> A_IWL<5710> A_IWL<5709> A_IWL<5708> A_IWL<5707> A_IWL<5706> A_IWL<5705> A_IWL<5704> A_IWL<5703> A_IWL<5702> A_IWL<5701> A_IWL<5700> A_IWL<5699> A_IWL<5698> A_IWL<5697> A_IWL<5696> A_IWL<5695> A_IWL<5694> A_IWL<5693> A_IWL<5692> A_IWL<5691> A_IWL<5690> A_IWL<5689> A_IWL<5688> A_IWL<5687> A_IWL<5686> A_IWL<5685> A_IWL<5684> A_IWL<5683> A_IWL<5682> A_IWL<5681> A_IWL<5680> A_IWL<5679> A_IWL<5678> A_IWL<5677> A_IWL<5676> A_IWL<5675> A_IWL<5674> A_IWL<5673> A_IWL<5672> A_IWL<5671> A_IWL<5670> A_IWL<5669> A_IWL<5668> A_IWL<5667> A_IWL<5666> A_IWL<5665> A_IWL<5664> A_IWL<5663> A_IWL<5662> A_IWL<5661> A_IWL<5660> A_IWL<5659> A_IWL<5658> A_IWL<5657> A_IWL<5656> A_IWL<5655> A_IWL<5654> A_IWL<5653> A_IWL<5652> A_IWL<5651> A_IWL<5650> A_IWL<5649> A_IWL<5648> A_IWL<5647> A_IWL<5646> A_IWL<5645> A_IWL<5644> A_IWL<5643> A_IWL<5642> A_IWL<5641> A_IWL<5640> A_IWL<5639> A_IWL<5638> A_IWL<5637> A_IWL<5636> A_IWL<5635> A_IWL<5634> A_IWL<5633> A_IWL<5632> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<21> A_BLC<43> A_BLC<42> A_BLC_TOP<43> A_BLC_TOP<42> A_BLT<43> A_BLT<42> A_BLT_TOP<43> A_BLT_TOP<42> A_IWL<5375> A_IWL<5374> A_IWL<5373> A_IWL<5372> A_IWL<5371> A_IWL<5370> A_IWL<5369> A_IWL<5368> A_IWL<5367> A_IWL<5366> A_IWL<5365> A_IWL<5364> A_IWL<5363> A_IWL<5362> A_IWL<5361> A_IWL<5360> A_IWL<5359> A_IWL<5358> A_IWL<5357> A_IWL<5356> A_IWL<5355> A_IWL<5354> A_IWL<5353> A_IWL<5352> A_IWL<5351> A_IWL<5350> A_IWL<5349> A_IWL<5348> A_IWL<5347> A_IWL<5346> A_IWL<5345> A_IWL<5344> A_IWL<5343> A_IWL<5342> A_IWL<5341> A_IWL<5340> A_IWL<5339> A_IWL<5338> A_IWL<5337> A_IWL<5336> A_IWL<5335> A_IWL<5334> A_IWL<5333> A_IWL<5332> A_IWL<5331> A_IWL<5330> A_IWL<5329> A_IWL<5328> A_IWL<5327> A_IWL<5326> A_IWL<5325> A_IWL<5324> A_IWL<5323> A_IWL<5322> A_IWL<5321> A_IWL<5320> A_IWL<5319> A_IWL<5318> A_IWL<5317> A_IWL<5316> A_IWL<5315> A_IWL<5314> A_IWL<5313> A_IWL<5312> A_IWL<5311> A_IWL<5310> A_IWL<5309> A_IWL<5308> A_IWL<5307> A_IWL<5306> A_IWL<5305> A_IWL<5304> A_IWL<5303> A_IWL<5302> A_IWL<5301> A_IWL<5300> A_IWL<5299> A_IWL<5298> A_IWL<5297> A_IWL<5296> A_IWL<5295> A_IWL<5294> A_IWL<5293> A_IWL<5292> A_IWL<5291> A_IWL<5290> A_IWL<5289> A_IWL<5288> A_IWL<5287> A_IWL<5286> A_IWL<5285> A_IWL<5284> A_IWL<5283> A_IWL<5282> A_IWL<5281> A_IWL<5280> A_IWL<5279> A_IWL<5278> A_IWL<5277> A_IWL<5276> A_IWL<5275> A_IWL<5274> A_IWL<5273> A_IWL<5272> A_IWL<5271> A_IWL<5270> A_IWL<5269> A_IWL<5268> A_IWL<5267> A_IWL<5266> A_IWL<5265> A_IWL<5264> A_IWL<5263> A_IWL<5262> A_IWL<5261> A_IWL<5260> A_IWL<5259> A_IWL<5258> A_IWL<5257> A_IWL<5256> A_IWL<5255> A_IWL<5254> A_IWL<5253> A_IWL<5252> A_IWL<5251> A_IWL<5250> A_IWL<5249> A_IWL<5248> A_IWL<5247> A_IWL<5246> A_IWL<5245> A_IWL<5244> A_IWL<5243> A_IWL<5242> A_IWL<5241> A_IWL<5240> A_IWL<5239> A_IWL<5238> A_IWL<5237> A_IWL<5236> A_IWL<5235> A_IWL<5234> A_IWL<5233> A_IWL<5232> A_IWL<5231> A_IWL<5230> A_IWL<5229> A_IWL<5228> A_IWL<5227> A_IWL<5226> A_IWL<5225> A_IWL<5224> A_IWL<5223> A_IWL<5222> A_IWL<5221> A_IWL<5220> A_IWL<5219> A_IWL<5218> A_IWL<5217> A_IWL<5216> A_IWL<5215> A_IWL<5214> A_IWL<5213> A_IWL<5212> A_IWL<5211> A_IWL<5210> A_IWL<5209> A_IWL<5208> A_IWL<5207> A_IWL<5206> A_IWL<5205> A_IWL<5204> A_IWL<5203> A_IWL<5202> A_IWL<5201> A_IWL<5200> A_IWL<5199> A_IWL<5198> A_IWL<5197> A_IWL<5196> A_IWL<5195> A_IWL<5194> A_IWL<5193> A_IWL<5192> A_IWL<5191> A_IWL<5190> A_IWL<5189> A_IWL<5188> A_IWL<5187> A_IWL<5186> A_IWL<5185> A_IWL<5184> A_IWL<5183> A_IWL<5182> A_IWL<5181> A_IWL<5180> A_IWL<5179> A_IWL<5178> A_IWL<5177> A_IWL<5176> A_IWL<5175> A_IWL<5174> A_IWL<5173> A_IWL<5172> A_IWL<5171> A_IWL<5170> A_IWL<5169> A_IWL<5168> A_IWL<5167> A_IWL<5166> A_IWL<5165> A_IWL<5164> A_IWL<5163> A_IWL<5162> A_IWL<5161> A_IWL<5160> A_IWL<5159> A_IWL<5158> A_IWL<5157> A_IWL<5156> A_IWL<5155> A_IWL<5154> A_IWL<5153> A_IWL<5152> A_IWL<5151> A_IWL<5150> A_IWL<5149> A_IWL<5148> A_IWL<5147> A_IWL<5146> A_IWL<5145> A_IWL<5144> A_IWL<5143> A_IWL<5142> A_IWL<5141> A_IWL<5140> A_IWL<5139> A_IWL<5138> A_IWL<5137> A_IWL<5136> A_IWL<5135> A_IWL<5134> A_IWL<5133> A_IWL<5132> A_IWL<5131> A_IWL<5130> A_IWL<5129> A_IWL<5128> A_IWL<5127> A_IWL<5126> A_IWL<5125> A_IWL<5124> A_IWL<5123> A_IWL<5122> A_IWL<5121> A_IWL<5120> A_IWL<5631> A_IWL<5630> A_IWL<5629> A_IWL<5628> A_IWL<5627> A_IWL<5626> A_IWL<5625> A_IWL<5624> A_IWL<5623> A_IWL<5622> A_IWL<5621> A_IWL<5620> A_IWL<5619> A_IWL<5618> A_IWL<5617> A_IWL<5616> A_IWL<5615> A_IWL<5614> A_IWL<5613> A_IWL<5612> A_IWL<5611> A_IWL<5610> A_IWL<5609> A_IWL<5608> A_IWL<5607> A_IWL<5606> A_IWL<5605> A_IWL<5604> A_IWL<5603> A_IWL<5602> A_IWL<5601> A_IWL<5600> A_IWL<5599> A_IWL<5598> A_IWL<5597> A_IWL<5596> A_IWL<5595> A_IWL<5594> A_IWL<5593> A_IWL<5592> A_IWL<5591> A_IWL<5590> A_IWL<5589> A_IWL<5588> A_IWL<5587> A_IWL<5586> A_IWL<5585> A_IWL<5584> A_IWL<5583> A_IWL<5582> A_IWL<5581> A_IWL<5580> A_IWL<5579> A_IWL<5578> A_IWL<5577> A_IWL<5576> A_IWL<5575> A_IWL<5574> A_IWL<5573> A_IWL<5572> A_IWL<5571> A_IWL<5570> A_IWL<5569> A_IWL<5568> A_IWL<5567> A_IWL<5566> A_IWL<5565> A_IWL<5564> A_IWL<5563> A_IWL<5562> A_IWL<5561> A_IWL<5560> A_IWL<5559> A_IWL<5558> A_IWL<5557> A_IWL<5556> A_IWL<5555> A_IWL<5554> A_IWL<5553> A_IWL<5552> A_IWL<5551> A_IWL<5550> A_IWL<5549> A_IWL<5548> A_IWL<5547> A_IWL<5546> A_IWL<5545> A_IWL<5544> A_IWL<5543> A_IWL<5542> A_IWL<5541> A_IWL<5540> A_IWL<5539> A_IWL<5538> A_IWL<5537> A_IWL<5536> A_IWL<5535> A_IWL<5534> A_IWL<5533> A_IWL<5532> A_IWL<5531> A_IWL<5530> A_IWL<5529> A_IWL<5528> A_IWL<5527> A_IWL<5526> A_IWL<5525> A_IWL<5524> A_IWL<5523> A_IWL<5522> A_IWL<5521> A_IWL<5520> A_IWL<5519> A_IWL<5518> A_IWL<5517> A_IWL<5516> A_IWL<5515> A_IWL<5514> A_IWL<5513> A_IWL<5512> A_IWL<5511> A_IWL<5510> A_IWL<5509> A_IWL<5508> A_IWL<5507> A_IWL<5506> A_IWL<5505> A_IWL<5504> A_IWL<5503> A_IWL<5502> A_IWL<5501> A_IWL<5500> A_IWL<5499> A_IWL<5498> A_IWL<5497> A_IWL<5496> A_IWL<5495> A_IWL<5494> A_IWL<5493> A_IWL<5492> A_IWL<5491> A_IWL<5490> A_IWL<5489> A_IWL<5488> A_IWL<5487> A_IWL<5486> A_IWL<5485> A_IWL<5484> A_IWL<5483> A_IWL<5482> A_IWL<5481> A_IWL<5480> A_IWL<5479> A_IWL<5478> A_IWL<5477> A_IWL<5476> A_IWL<5475> A_IWL<5474> A_IWL<5473> A_IWL<5472> A_IWL<5471> A_IWL<5470> A_IWL<5469> A_IWL<5468> A_IWL<5467> A_IWL<5466> A_IWL<5465> A_IWL<5464> A_IWL<5463> A_IWL<5462> A_IWL<5461> A_IWL<5460> A_IWL<5459> A_IWL<5458> A_IWL<5457> A_IWL<5456> A_IWL<5455> A_IWL<5454> A_IWL<5453> A_IWL<5452> A_IWL<5451> A_IWL<5450> A_IWL<5449> A_IWL<5448> A_IWL<5447> A_IWL<5446> A_IWL<5445> A_IWL<5444> A_IWL<5443> A_IWL<5442> A_IWL<5441> A_IWL<5440> A_IWL<5439> A_IWL<5438> A_IWL<5437> A_IWL<5436> A_IWL<5435> A_IWL<5434> A_IWL<5433> A_IWL<5432> A_IWL<5431> A_IWL<5430> A_IWL<5429> A_IWL<5428> A_IWL<5427> A_IWL<5426> A_IWL<5425> A_IWL<5424> A_IWL<5423> A_IWL<5422> A_IWL<5421> A_IWL<5420> A_IWL<5419> A_IWL<5418> A_IWL<5417> A_IWL<5416> A_IWL<5415> A_IWL<5414> A_IWL<5413> A_IWL<5412> A_IWL<5411> A_IWL<5410> A_IWL<5409> A_IWL<5408> A_IWL<5407> A_IWL<5406> A_IWL<5405> A_IWL<5404> A_IWL<5403> A_IWL<5402> A_IWL<5401> A_IWL<5400> A_IWL<5399> A_IWL<5398> A_IWL<5397> A_IWL<5396> A_IWL<5395> A_IWL<5394> A_IWL<5393> A_IWL<5392> A_IWL<5391> A_IWL<5390> A_IWL<5389> A_IWL<5388> A_IWL<5387> A_IWL<5386> A_IWL<5385> A_IWL<5384> A_IWL<5383> A_IWL<5382> A_IWL<5381> A_IWL<5380> A_IWL<5379> A_IWL<5378> A_IWL<5377> A_IWL<5376> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<20> A_BLC<41> A_BLC<40> A_BLC_TOP<41> A_BLC_TOP<40> A_BLT<41> A_BLT<40> A_BLT_TOP<41> A_BLT_TOP<40> A_IWL<5119> A_IWL<5118> A_IWL<5117> A_IWL<5116> A_IWL<5115> A_IWL<5114> A_IWL<5113> A_IWL<5112> A_IWL<5111> A_IWL<5110> A_IWL<5109> A_IWL<5108> A_IWL<5107> A_IWL<5106> A_IWL<5105> A_IWL<5104> A_IWL<5103> A_IWL<5102> A_IWL<5101> A_IWL<5100> A_IWL<5099> A_IWL<5098> A_IWL<5097> A_IWL<5096> A_IWL<5095> A_IWL<5094> A_IWL<5093> A_IWL<5092> A_IWL<5091> A_IWL<5090> A_IWL<5089> A_IWL<5088> A_IWL<5087> A_IWL<5086> A_IWL<5085> A_IWL<5084> A_IWL<5083> A_IWL<5082> A_IWL<5081> A_IWL<5080> A_IWL<5079> A_IWL<5078> A_IWL<5077> A_IWL<5076> A_IWL<5075> A_IWL<5074> A_IWL<5073> A_IWL<5072> A_IWL<5071> A_IWL<5070> A_IWL<5069> A_IWL<5068> A_IWL<5067> A_IWL<5066> A_IWL<5065> A_IWL<5064> A_IWL<5063> A_IWL<5062> A_IWL<5061> A_IWL<5060> A_IWL<5059> A_IWL<5058> A_IWL<5057> A_IWL<5056> A_IWL<5055> A_IWL<5054> A_IWL<5053> A_IWL<5052> A_IWL<5051> A_IWL<5050> A_IWL<5049> A_IWL<5048> A_IWL<5047> A_IWL<5046> A_IWL<5045> A_IWL<5044> A_IWL<5043> A_IWL<5042> A_IWL<5041> A_IWL<5040> A_IWL<5039> A_IWL<5038> A_IWL<5037> A_IWL<5036> A_IWL<5035> A_IWL<5034> A_IWL<5033> A_IWL<5032> A_IWL<5031> A_IWL<5030> A_IWL<5029> A_IWL<5028> A_IWL<5027> A_IWL<5026> A_IWL<5025> A_IWL<5024> A_IWL<5023> A_IWL<5022> A_IWL<5021> A_IWL<5020> A_IWL<5019> A_IWL<5018> A_IWL<5017> A_IWL<5016> A_IWL<5015> A_IWL<5014> A_IWL<5013> A_IWL<5012> A_IWL<5011> A_IWL<5010> A_IWL<5009> A_IWL<5008> A_IWL<5007> A_IWL<5006> A_IWL<5005> A_IWL<5004> A_IWL<5003> A_IWL<5002> A_IWL<5001> A_IWL<5000> A_IWL<4999> A_IWL<4998> A_IWL<4997> A_IWL<4996> A_IWL<4995> A_IWL<4994> A_IWL<4993> A_IWL<4992> A_IWL<4991> A_IWL<4990> A_IWL<4989> A_IWL<4988> A_IWL<4987> A_IWL<4986> A_IWL<4985> A_IWL<4984> A_IWL<4983> A_IWL<4982> A_IWL<4981> A_IWL<4980> A_IWL<4979> A_IWL<4978> A_IWL<4977> A_IWL<4976> A_IWL<4975> A_IWL<4974> A_IWL<4973> A_IWL<4972> A_IWL<4971> A_IWL<4970> A_IWL<4969> A_IWL<4968> A_IWL<4967> A_IWL<4966> A_IWL<4965> A_IWL<4964> A_IWL<4963> A_IWL<4962> A_IWL<4961> A_IWL<4960> A_IWL<4959> A_IWL<4958> A_IWL<4957> A_IWL<4956> A_IWL<4955> A_IWL<4954> A_IWL<4953> A_IWL<4952> A_IWL<4951> A_IWL<4950> A_IWL<4949> A_IWL<4948> A_IWL<4947> A_IWL<4946> A_IWL<4945> A_IWL<4944> A_IWL<4943> A_IWL<4942> A_IWL<4941> A_IWL<4940> A_IWL<4939> A_IWL<4938> A_IWL<4937> A_IWL<4936> A_IWL<4935> A_IWL<4934> A_IWL<4933> A_IWL<4932> A_IWL<4931> A_IWL<4930> A_IWL<4929> A_IWL<4928> A_IWL<4927> A_IWL<4926> A_IWL<4925> A_IWL<4924> A_IWL<4923> A_IWL<4922> A_IWL<4921> A_IWL<4920> A_IWL<4919> A_IWL<4918> A_IWL<4917> A_IWL<4916> A_IWL<4915> A_IWL<4914> A_IWL<4913> A_IWL<4912> A_IWL<4911> A_IWL<4910> A_IWL<4909> A_IWL<4908> A_IWL<4907> A_IWL<4906> A_IWL<4905> A_IWL<4904> A_IWL<4903> A_IWL<4902> A_IWL<4901> A_IWL<4900> A_IWL<4899> A_IWL<4898> A_IWL<4897> A_IWL<4896> A_IWL<4895> A_IWL<4894> A_IWL<4893> A_IWL<4892> A_IWL<4891> A_IWL<4890> A_IWL<4889> A_IWL<4888> A_IWL<4887> A_IWL<4886> A_IWL<4885> A_IWL<4884> A_IWL<4883> A_IWL<4882> A_IWL<4881> A_IWL<4880> A_IWL<4879> A_IWL<4878> A_IWL<4877> A_IWL<4876> A_IWL<4875> A_IWL<4874> A_IWL<4873> A_IWL<4872> A_IWL<4871> A_IWL<4870> A_IWL<4869> A_IWL<4868> A_IWL<4867> A_IWL<4866> A_IWL<4865> A_IWL<4864> A_IWL<5375> A_IWL<5374> A_IWL<5373> A_IWL<5372> A_IWL<5371> A_IWL<5370> A_IWL<5369> A_IWL<5368> A_IWL<5367> A_IWL<5366> A_IWL<5365> A_IWL<5364> A_IWL<5363> A_IWL<5362> A_IWL<5361> A_IWL<5360> A_IWL<5359> A_IWL<5358> A_IWL<5357> A_IWL<5356> A_IWL<5355> A_IWL<5354> A_IWL<5353> A_IWL<5352> A_IWL<5351> A_IWL<5350> A_IWL<5349> A_IWL<5348> A_IWL<5347> A_IWL<5346> A_IWL<5345> A_IWL<5344> A_IWL<5343> A_IWL<5342> A_IWL<5341> A_IWL<5340> A_IWL<5339> A_IWL<5338> A_IWL<5337> A_IWL<5336> A_IWL<5335> A_IWL<5334> A_IWL<5333> A_IWL<5332> A_IWL<5331> A_IWL<5330> A_IWL<5329> A_IWL<5328> A_IWL<5327> A_IWL<5326> A_IWL<5325> A_IWL<5324> A_IWL<5323> A_IWL<5322> A_IWL<5321> A_IWL<5320> A_IWL<5319> A_IWL<5318> A_IWL<5317> A_IWL<5316> A_IWL<5315> A_IWL<5314> A_IWL<5313> A_IWL<5312> A_IWL<5311> A_IWL<5310> A_IWL<5309> A_IWL<5308> A_IWL<5307> A_IWL<5306> A_IWL<5305> A_IWL<5304> A_IWL<5303> A_IWL<5302> A_IWL<5301> A_IWL<5300> A_IWL<5299> A_IWL<5298> A_IWL<5297> A_IWL<5296> A_IWL<5295> A_IWL<5294> A_IWL<5293> A_IWL<5292> A_IWL<5291> A_IWL<5290> A_IWL<5289> A_IWL<5288> A_IWL<5287> A_IWL<5286> A_IWL<5285> A_IWL<5284> A_IWL<5283> A_IWL<5282> A_IWL<5281> A_IWL<5280> A_IWL<5279> A_IWL<5278> A_IWL<5277> A_IWL<5276> A_IWL<5275> A_IWL<5274> A_IWL<5273> A_IWL<5272> A_IWL<5271> A_IWL<5270> A_IWL<5269> A_IWL<5268> A_IWL<5267> A_IWL<5266> A_IWL<5265> A_IWL<5264> A_IWL<5263> A_IWL<5262> A_IWL<5261> A_IWL<5260> A_IWL<5259> A_IWL<5258> A_IWL<5257> A_IWL<5256> A_IWL<5255> A_IWL<5254> A_IWL<5253> A_IWL<5252> A_IWL<5251> A_IWL<5250> A_IWL<5249> A_IWL<5248> A_IWL<5247> A_IWL<5246> A_IWL<5245> A_IWL<5244> A_IWL<5243> A_IWL<5242> A_IWL<5241> A_IWL<5240> A_IWL<5239> A_IWL<5238> A_IWL<5237> A_IWL<5236> A_IWL<5235> A_IWL<5234> A_IWL<5233> A_IWL<5232> A_IWL<5231> A_IWL<5230> A_IWL<5229> A_IWL<5228> A_IWL<5227> A_IWL<5226> A_IWL<5225> A_IWL<5224> A_IWL<5223> A_IWL<5222> A_IWL<5221> A_IWL<5220> A_IWL<5219> A_IWL<5218> A_IWL<5217> A_IWL<5216> A_IWL<5215> A_IWL<5214> A_IWL<5213> A_IWL<5212> A_IWL<5211> A_IWL<5210> A_IWL<5209> A_IWL<5208> A_IWL<5207> A_IWL<5206> A_IWL<5205> A_IWL<5204> A_IWL<5203> A_IWL<5202> A_IWL<5201> A_IWL<5200> A_IWL<5199> A_IWL<5198> A_IWL<5197> A_IWL<5196> A_IWL<5195> A_IWL<5194> A_IWL<5193> A_IWL<5192> A_IWL<5191> A_IWL<5190> A_IWL<5189> A_IWL<5188> A_IWL<5187> A_IWL<5186> A_IWL<5185> A_IWL<5184> A_IWL<5183> A_IWL<5182> A_IWL<5181> A_IWL<5180> A_IWL<5179> A_IWL<5178> A_IWL<5177> A_IWL<5176> A_IWL<5175> A_IWL<5174> A_IWL<5173> A_IWL<5172> A_IWL<5171> A_IWL<5170> A_IWL<5169> A_IWL<5168> A_IWL<5167> A_IWL<5166> A_IWL<5165> A_IWL<5164> A_IWL<5163> A_IWL<5162> A_IWL<5161> A_IWL<5160> A_IWL<5159> A_IWL<5158> A_IWL<5157> A_IWL<5156> A_IWL<5155> A_IWL<5154> A_IWL<5153> A_IWL<5152> A_IWL<5151> A_IWL<5150> A_IWL<5149> A_IWL<5148> A_IWL<5147> A_IWL<5146> A_IWL<5145> A_IWL<5144> A_IWL<5143> A_IWL<5142> A_IWL<5141> A_IWL<5140> A_IWL<5139> A_IWL<5138> A_IWL<5137> A_IWL<5136> A_IWL<5135> A_IWL<5134> A_IWL<5133> A_IWL<5132> A_IWL<5131> A_IWL<5130> A_IWL<5129> A_IWL<5128> A_IWL<5127> A_IWL<5126> A_IWL<5125> A_IWL<5124> A_IWL<5123> A_IWL<5122> A_IWL<5121> A_IWL<5120> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<19> A_BLC<39> A_BLC<38> A_BLC_TOP<39> A_BLC_TOP<38> A_BLT<39> A_BLT<38> A_BLT_TOP<39> A_BLT_TOP<38> A_IWL<4863> A_IWL<4862> A_IWL<4861> A_IWL<4860> A_IWL<4859> A_IWL<4858> A_IWL<4857> A_IWL<4856> A_IWL<4855> A_IWL<4854> A_IWL<4853> A_IWL<4852> A_IWL<4851> A_IWL<4850> A_IWL<4849> A_IWL<4848> A_IWL<4847> A_IWL<4846> A_IWL<4845> A_IWL<4844> A_IWL<4843> A_IWL<4842> A_IWL<4841> A_IWL<4840> A_IWL<4839> A_IWL<4838> A_IWL<4837> A_IWL<4836> A_IWL<4835> A_IWL<4834> A_IWL<4833> A_IWL<4832> A_IWL<4831> A_IWL<4830> A_IWL<4829> A_IWL<4828> A_IWL<4827> A_IWL<4826> A_IWL<4825> A_IWL<4824> A_IWL<4823> A_IWL<4822> A_IWL<4821> A_IWL<4820> A_IWL<4819> A_IWL<4818> A_IWL<4817> A_IWL<4816> A_IWL<4815> A_IWL<4814> A_IWL<4813> A_IWL<4812> A_IWL<4811> A_IWL<4810> A_IWL<4809> A_IWL<4808> A_IWL<4807> A_IWL<4806> A_IWL<4805> A_IWL<4804> A_IWL<4803> A_IWL<4802> A_IWL<4801> A_IWL<4800> A_IWL<4799> A_IWL<4798> A_IWL<4797> A_IWL<4796> A_IWL<4795> A_IWL<4794> A_IWL<4793> A_IWL<4792> A_IWL<4791> A_IWL<4790> A_IWL<4789> A_IWL<4788> A_IWL<4787> A_IWL<4786> A_IWL<4785> A_IWL<4784> A_IWL<4783> A_IWL<4782> A_IWL<4781> A_IWL<4780> A_IWL<4779> A_IWL<4778> A_IWL<4777> A_IWL<4776> A_IWL<4775> A_IWL<4774> A_IWL<4773> A_IWL<4772> A_IWL<4771> A_IWL<4770> A_IWL<4769> A_IWL<4768> A_IWL<4767> A_IWL<4766> A_IWL<4765> A_IWL<4764> A_IWL<4763> A_IWL<4762> A_IWL<4761> A_IWL<4760> A_IWL<4759> A_IWL<4758> A_IWL<4757> A_IWL<4756> A_IWL<4755> A_IWL<4754> A_IWL<4753> A_IWL<4752> A_IWL<4751> A_IWL<4750> A_IWL<4749> A_IWL<4748> A_IWL<4747> A_IWL<4746> A_IWL<4745> A_IWL<4744> A_IWL<4743> A_IWL<4742> A_IWL<4741> A_IWL<4740> A_IWL<4739> A_IWL<4738> A_IWL<4737> A_IWL<4736> A_IWL<4735> A_IWL<4734> A_IWL<4733> A_IWL<4732> A_IWL<4731> A_IWL<4730> A_IWL<4729> A_IWL<4728> A_IWL<4727> A_IWL<4726> A_IWL<4725> A_IWL<4724> A_IWL<4723> A_IWL<4722> A_IWL<4721> A_IWL<4720> A_IWL<4719> A_IWL<4718> A_IWL<4717> A_IWL<4716> A_IWL<4715> A_IWL<4714> A_IWL<4713> A_IWL<4712> A_IWL<4711> A_IWL<4710> A_IWL<4709> A_IWL<4708> A_IWL<4707> A_IWL<4706> A_IWL<4705> A_IWL<4704> A_IWL<4703> A_IWL<4702> A_IWL<4701> A_IWL<4700> A_IWL<4699> A_IWL<4698> A_IWL<4697> A_IWL<4696> A_IWL<4695> A_IWL<4694> A_IWL<4693> A_IWL<4692> A_IWL<4691> A_IWL<4690> A_IWL<4689> A_IWL<4688> A_IWL<4687> A_IWL<4686> A_IWL<4685> A_IWL<4684> A_IWL<4683> A_IWL<4682> A_IWL<4681> A_IWL<4680> A_IWL<4679> A_IWL<4678> A_IWL<4677> A_IWL<4676> A_IWL<4675> A_IWL<4674> A_IWL<4673> A_IWL<4672> A_IWL<4671> A_IWL<4670> A_IWL<4669> A_IWL<4668> A_IWL<4667> A_IWL<4666> A_IWL<4665> A_IWL<4664> A_IWL<4663> A_IWL<4662> A_IWL<4661> A_IWL<4660> A_IWL<4659> A_IWL<4658> A_IWL<4657> A_IWL<4656> A_IWL<4655> A_IWL<4654> A_IWL<4653> A_IWL<4652> A_IWL<4651> A_IWL<4650> A_IWL<4649> A_IWL<4648> A_IWL<4647> A_IWL<4646> A_IWL<4645> A_IWL<4644> A_IWL<4643> A_IWL<4642> A_IWL<4641> A_IWL<4640> A_IWL<4639> A_IWL<4638> A_IWL<4637> A_IWL<4636> A_IWL<4635> A_IWL<4634> A_IWL<4633> A_IWL<4632> A_IWL<4631> A_IWL<4630> A_IWL<4629> A_IWL<4628> A_IWL<4627> A_IWL<4626> A_IWL<4625> A_IWL<4624> A_IWL<4623> A_IWL<4622> A_IWL<4621> A_IWL<4620> A_IWL<4619> A_IWL<4618> A_IWL<4617> A_IWL<4616> A_IWL<4615> A_IWL<4614> A_IWL<4613> A_IWL<4612> A_IWL<4611> A_IWL<4610> A_IWL<4609> A_IWL<4608> A_IWL<5119> A_IWL<5118> A_IWL<5117> A_IWL<5116> A_IWL<5115> A_IWL<5114> A_IWL<5113> A_IWL<5112> A_IWL<5111> A_IWL<5110> A_IWL<5109> A_IWL<5108> A_IWL<5107> A_IWL<5106> A_IWL<5105> A_IWL<5104> A_IWL<5103> A_IWL<5102> A_IWL<5101> A_IWL<5100> A_IWL<5099> A_IWL<5098> A_IWL<5097> A_IWL<5096> A_IWL<5095> A_IWL<5094> A_IWL<5093> A_IWL<5092> A_IWL<5091> A_IWL<5090> A_IWL<5089> A_IWL<5088> A_IWL<5087> A_IWL<5086> A_IWL<5085> A_IWL<5084> A_IWL<5083> A_IWL<5082> A_IWL<5081> A_IWL<5080> A_IWL<5079> A_IWL<5078> A_IWL<5077> A_IWL<5076> A_IWL<5075> A_IWL<5074> A_IWL<5073> A_IWL<5072> A_IWL<5071> A_IWL<5070> A_IWL<5069> A_IWL<5068> A_IWL<5067> A_IWL<5066> A_IWL<5065> A_IWL<5064> A_IWL<5063> A_IWL<5062> A_IWL<5061> A_IWL<5060> A_IWL<5059> A_IWL<5058> A_IWL<5057> A_IWL<5056> A_IWL<5055> A_IWL<5054> A_IWL<5053> A_IWL<5052> A_IWL<5051> A_IWL<5050> A_IWL<5049> A_IWL<5048> A_IWL<5047> A_IWL<5046> A_IWL<5045> A_IWL<5044> A_IWL<5043> A_IWL<5042> A_IWL<5041> A_IWL<5040> A_IWL<5039> A_IWL<5038> A_IWL<5037> A_IWL<5036> A_IWL<5035> A_IWL<5034> A_IWL<5033> A_IWL<5032> A_IWL<5031> A_IWL<5030> A_IWL<5029> A_IWL<5028> A_IWL<5027> A_IWL<5026> A_IWL<5025> A_IWL<5024> A_IWL<5023> A_IWL<5022> A_IWL<5021> A_IWL<5020> A_IWL<5019> A_IWL<5018> A_IWL<5017> A_IWL<5016> A_IWL<5015> A_IWL<5014> A_IWL<5013> A_IWL<5012> A_IWL<5011> A_IWL<5010> A_IWL<5009> A_IWL<5008> A_IWL<5007> A_IWL<5006> A_IWL<5005> A_IWL<5004> A_IWL<5003> A_IWL<5002> A_IWL<5001> A_IWL<5000> A_IWL<4999> A_IWL<4998> A_IWL<4997> A_IWL<4996> A_IWL<4995> A_IWL<4994> A_IWL<4993> A_IWL<4992> A_IWL<4991> A_IWL<4990> A_IWL<4989> A_IWL<4988> A_IWL<4987> A_IWL<4986> A_IWL<4985> A_IWL<4984> A_IWL<4983> A_IWL<4982> A_IWL<4981> A_IWL<4980> A_IWL<4979> A_IWL<4978> A_IWL<4977> A_IWL<4976> A_IWL<4975> A_IWL<4974> A_IWL<4973> A_IWL<4972> A_IWL<4971> A_IWL<4970> A_IWL<4969> A_IWL<4968> A_IWL<4967> A_IWL<4966> A_IWL<4965> A_IWL<4964> A_IWL<4963> A_IWL<4962> A_IWL<4961> A_IWL<4960> A_IWL<4959> A_IWL<4958> A_IWL<4957> A_IWL<4956> A_IWL<4955> A_IWL<4954> A_IWL<4953> A_IWL<4952> A_IWL<4951> A_IWL<4950> A_IWL<4949> A_IWL<4948> A_IWL<4947> A_IWL<4946> A_IWL<4945> A_IWL<4944> A_IWL<4943> A_IWL<4942> A_IWL<4941> A_IWL<4940> A_IWL<4939> A_IWL<4938> A_IWL<4937> A_IWL<4936> A_IWL<4935> A_IWL<4934> A_IWL<4933> A_IWL<4932> A_IWL<4931> A_IWL<4930> A_IWL<4929> A_IWL<4928> A_IWL<4927> A_IWL<4926> A_IWL<4925> A_IWL<4924> A_IWL<4923> A_IWL<4922> A_IWL<4921> A_IWL<4920> A_IWL<4919> A_IWL<4918> A_IWL<4917> A_IWL<4916> A_IWL<4915> A_IWL<4914> A_IWL<4913> A_IWL<4912> A_IWL<4911> A_IWL<4910> A_IWL<4909> A_IWL<4908> A_IWL<4907> A_IWL<4906> A_IWL<4905> A_IWL<4904> A_IWL<4903> A_IWL<4902> A_IWL<4901> A_IWL<4900> A_IWL<4899> A_IWL<4898> A_IWL<4897> A_IWL<4896> A_IWL<4895> A_IWL<4894> A_IWL<4893> A_IWL<4892> A_IWL<4891> A_IWL<4890> A_IWL<4889> A_IWL<4888> A_IWL<4887> A_IWL<4886> A_IWL<4885> A_IWL<4884> A_IWL<4883> A_IWL<4882> A_IWL<4881> A_IWL<4880> A_IWL<4879> A_IWL<4878> A_IWL<4877> A_IWL<4876> A_IWL<4875> A_IWL<4874> A_IWL<4873> A_IWL<4872> A_IWL<4871> A_IWL<4870> A_IWL<4869> A_IWL<4868> A_IWL<4867> A_IWL<4866> A_IWL<4865> A_IWL<4864> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<18> A_BLC<37> A_BLC<36> A_BLC_TOP<37> A_BLC_TOP<36> A_BLT<37> A_BLT<36> A_BLT_TOP<37> A_BLT_TOP<36> A_IWL<4607> A_IWL<4606> A_IWL<4605> A_IWL<4604> A_IWL<4603> A_IWL<4602> A_IWL<4601> A_IWL<4600> A_IWL<4599> A_IWL<4598> A_IWL<4597> A_IWL<4596> A_IWL<4595> A_IWL<4594> A_IWL<4593> A_IWL<4592> A_IWL<4591> A_IWL<4590> A_IWL<4589> A_IWL<4588> A_IWL<4587> A_IWL<4586> A_IWL<4585> A_IWL<4584> A_IWL<4583> A_IWL<4582> A_IWL<4581> A_IWL<4580> A_IWL<4579> A_IWL<4578> A_IWL<4577> A_IWL<4576> A_IWL<4575> A_IWL<4574> A_IWL<4573> A_IWL<4572> A_IWL<4571> A_IWL<4570> A_IWL<4569> A_IWL<4568> A_IWL<4567> A_IWL<4566> A_IWL<4565> A_IWL<4564> A_IWL<4563> A_IWL<4562> A_IWL<4561> A_IWL<4560> A_IWL<4559> A_IWL<4558> A_IWL<4557> A_IWL<4556> A_IWL<4555> A_IWL<4554> A_IWL<4553> A_IWL<4552> A_IWL<4551> A_IWL<4550> A_IWL<4549> A_IWL<4548> A_IWL<4547> A_IWL<4546> A_IWL<4545> A_IWL<4544> A_IWL<4543> A_IWL<4542> A_IWL<4541> A_IWL<4540> A_IWL<4539> A_IWL<4538> A_IWL<4537> A_IWL<4536> A_IWL<4535> A_IWL<4534> A_IWL<4533> A_IWL<4532> A_IWL<4531> A_IWL<4530> A_IWL<4529> A_IWL<4528> A_IWL<4527> A_IWL<4526> A_IWL<4525> A_IWL<4524> A_IWL<4523> A_IWL<4522> A_IWL<4521> A_IWL<4520> A_IWL<4519> A_IWL<4518> A_IWL<4517> A_IWL<4516> A_IWL<4515> A_IWL<4514> A_IWL<4513> A_IWL<4512> A_IWL<4511> A_IWL<4510> A_IWL<4509> A_IWL<4508> A_IWL<4507> A_IWL<4506> A_IWL<4505> A_IWL<4504> A_IWL<4503> A_IWL<4502> A_IWL<4501> A_IWL<4500> A_IWL<4499> A_IWL<4498> A_IWL<4497> A_IWL<4496> A_IWL<4495> A_IWL<4494> A_IWL<4493> A_IWL<4492> A_IWL<4491> A_IWL<4490> A_IWL<4489> A_IWL<4488> A_IWL<4487> A_IWL<4486> A_IWL<4485> A_IWL<4484> A_IWL<4483> A_IWL<4482> A_IWL<4481> A_IWL<4480> A_IWL<4479> A_IWL<4478> A_IWL<4477> A_IWL<4476> A_IWL<4475> A_IWL<4474> A_IWL<4473> A_IWL<4472> A_IWL<4471> A_IWL<4470> A_IWL<4469> A_IWL<4468> A_IWL<4467> A_IWL<4466> A_IWL<4465> A_IWL<4464> A_IWL<4463> A_IWL<4462> A_IWL<4461> A_IWL<4460> A_IWL<4459> A_IWL<4458> A_IWL<4457> A_IWL<4456> A_IWL<4455> A_IWL<4454> A_IWL<4453> A_IWL<4452> A_IWL<4451> A_IWL<4450> A_IWL<4449> A_IWL<4448> A_IWL<4447> A_IWL<4446> A_IWL<4445> A_IWL<4444> A_IWL<4443> A_IWL<4442> A_IWL<4441> A_IWL<4440> A_IWL<4439> A_IWL<4438> A_IWL<4437> A_IWL<4436> A_IWL<4435> A_IWL<4434> A_IWL<4433> A_IWL<4432> A_IWL<4431> A_IWL<4430> A_IWL<4429> A_IWL<4428> A_IWL<4427> A_IWL<4426> A_IWL<4425> A_IWL<4424> A_IWL<4423> A_IWL<4422> A_IWL<4421> A_IWL<4420> A_IWL<4419> A_IWL<4418> A_IWL<4417> A_IWL<4416> A_IWL<4415> A_IWL<4414> A_IWL<4413> A_IWL<4412> A_IWL<4411> A_IWL<4410> A_IWL<4409> A_IWL<4408> A_IWL<4407> A_IWL<4406> A_IWL<4405> A_IWL<4404> A_IWL<4403> A_IWL<4402> A_IWL<4401> A_IWL<4400> A_IWL<4399> A_IWL<4398> A_IWL<4397> A_IWL<4396> A_IWL<4395> A_IWL<4394> A_IWL<4393> A_IWL<4392> A_IWL<4391> A_IWL<4390> A_IWL<4389> A_IWL<4388> A_IWL<4387> A_IWL<4386> A_IWL<4385> A_IWL<4384> A_IWL<4383> A_IWL<4382> A_IWL<4381> A_IWL<4380> A_IWL<4379> A_IWL<4378> A_IWL<4377> A_IWL<4376> A_IWL<4375> A_IWL<4374> A_IWL<4373> A_IWL<4372> A_IWL<4371> A_IWL<4370> A_IWL<4369> A_IWL<4368> A_IWL<4367> A_IWL<4366> A_IWL<4365> A_IWL<4364> A_IWL<4363> A_IWL<4362> A_IWL<4361> A_IWL<4360> A_IWL<4359> A_IWL<4358> A_IWL<4357> A_IWL<4356> A_IWL<4355> A_IWL<4354> A_IWL<4353> A_IWL<4352> A_IWL<4863> A_IWL<4862> A_IWL<4861> A_IWL<4860> A_IWL<4859> A_IWL<4858> A_IWL<4857> A_IWL<4856> A_IWL<4855> A_IWL<4854> A_IWL<4853> A_IWL<4852> A_IWL<4851> A_IWL<4850> A_IWL<4849> A_IWL<4848> A_IWL<4847> A_IWL<4846> A_IWL<4845> A_IWL<4844> A_IWL<4843> A_IWL<4842> A_IWL<4841> A_IWL<4840> A_IWL<4839> A_IWL<4838> A_IWL<4837> A_IWL<4836> A_IWL<4835> A_IWL<4834> A_IWL<4833> A_IWL<4832> A_IWL<4831> A_IWL<4830> A_IWL<4829> A_IWL<4828> A_IWL<4827> A_IWL<4826> A_IWL<4825> A_IWL<4824> A_IWL<4823> A_IWL<4822> A_IWL<4821> A_IWL<4820> A_IWL<4819> A_IWL<4818> A_IWL<4817> A_IWL<4816> A_IWL<4815> A_IWL<4814> A_IWL<4813> A_IWL<4812> A_IWL<4811> A_IWL<4810> A_IWL<4809> A_IWL<4808> A_IWL<4807> A_IWL<4806> A_IWL<4805> A_IWL<4804> A_IWL<4803> A_IWL<4802> A_IWL<4801> A_IWL<4800> A_IWL<4799> A_IWL<4798> A_IWL<4797> A_IWL<4796> A_IWL<4795> A_IWL<4794> A_IWL<4793> A_IWL<4792> A_IWL<4791> A_IWL<4790> A_IWL<4789> A_IWL<4788> A_IWL<4787> A_IWL<4786> A_IWL<4785> A_IWL<4784> A_IWL<4783> A_IWL<4782> A_IWL<4781> A_IWL<4780> A_IWL<4779> A_IWL<4778> A_IWL<4777> A_IWL<4776> A_IWL<4775> A_IWL<4774> A_IWL<4773> A_IWL<4772> A_IWL<4771> A_IWL<4770> A_IWL<4769> A_IWL<4768> A_IWL<4767> A_IWL<4766> A_IWL<4765> A_IWL<4764> A_IWL<4763> A_IWL<4762> A_IWL<4761> A_IWL<4760> A_IWL<4759> A_IWL<4758> A_IWL<4757> A_IWL<4756> A_IWL<4755> A_IWL<4754> A_IWL<4753> A_IWL<4752> A_IWL<4751> A_IWL<4750> A_IWL<4749> A_IWL<4748> A_IWL<4747> A_IWL<4746> A_IWL<4745> A_IWL<4744> A_IWL<4743> A_IWL<4742> A_IWL<4741> A_IWL<4740> A_IWL<4739> A_IWL<4738> A_IWL<4737> A_IWL<4736> A_IWL<4735> A_IWL<4734> A_IWL<4733> A_IWL<4732> A_IWL<4731> A_IWL<4730> A_IWL<4729> A_IWL<4728> A_IWL<4727> A_IWL<4726> A_IWL<4725> A_IWL<4724> A_IWL<4723> A_IWL<4722> A_IWL<4721> A_IWL<4720> A_IWL<4719> A_IWL<4718> A_IWL<4717> A_IWL<4716> A_IWL<4715> A_IWL<4714> A_IWL<4713> A_IWL<4712> A_IWL<4711> A_IWL<4710> A_IWL<4709> A_IWL<4708> A_IWL<4707> A_IWL<4706> A_IWL<4705> A_IWL<4704> A_IWL<4703> A_IWL<4702> A_IWL<4701> A_IWL<4700> A_IWL<4699> A_IWL<4698> A_IWL<4697> A_IWL<4696> A_IWL<4695> A_IWL<4694> A_IWL<4693> A_IWL<4692> A_IWL<4691> A_IWL<4690> A_IWL<4689> A_IWL<4688> A_IWL<4687> A_IWL<4686> A_IWL<4685> A_IWL<4684> A_IWL<4683> A_IWL<4682> A_IWL<4681> A_IWL<4680> A_IWL<4679> A_IWL<4678> A_IWL<4677> A_IWL<4676> A_IWL<4675> A_IWL<4674> A_IWL<4673> A_IWL<4672> A_IWL<4671> A_IWL<4670> A_IWL<4669> A_IWL<4668> A_IWL<4667> A_IWL<4666> A_IWL<4665> A_IWL<4664> A_IWL<4663> A_IWL<4662> A_IWL<4661> A_IWL<4660> A_IWL<4659> A_IWL<4658> A_IWL<4657> A_IWL<4656> A_IWL<4655> A_IWL<4654> A_IWL<4653> A_IWL<4652> A_IWL<4651> A_IWL<4650> A_IWL<4649> A_IWL<4648> A_IWL<4647> A_IWL<4646> A_IWL<4645> A_IWL<4644> A_IWL<4643> A_IWL<4642> A_IWL<4641> A_IWL<4640> A_IWL<4639> A_IWL<4638> A_IWL<4637> A_IWL<4636> A_IWL<4635> A_IWL<4634> A_IWL<4633> A_IWL<4632> A_IWL<4631> A_IWL<4630> A_IWL<4629> A_IWL<4628> A_IWL<4627> A_IWL<4626> A_IWL<4625> A_IWL<4624> A_IWL<4623> A_IWL<4622> A_IWL<4621> A_IWL<4620> A_IWL<4619> A_IWL<4618> A_IWL<4617> A_IWL<4616> A_IWL<4615> A_IWL<4614> A_IWL<4613> A_IWL<4612> A_IWL<4611> A_IWL<4610> A_IWL<4609> A_IWL<4608> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<17> A_BLC<35> A_BLC<34> A_BLC_TOP<35> A_BLC_TOP<34> A_BLT<35> A_BLT<34> A_BLT_TOP<35> A_BLT_TOP<34> A_IWL<4351> A_IWL<4350> A_IWL<4349> A_IWL<4348> A_IWL<4347> A_IWL<4346> A_IWL<4345> A_IWL<4344> A_IWL<4343> A_IWL<4342> A_IWL<4341> A_IWL<4340> A_IWL<4339> A_IWL<4338> A_IWL<4337> A_IWL<4336> A_IWL<4335> A_IWL<4334> A_IWL<4333> A_IWL<4332> A_IWL<4331> A_IWL<4330> A_IWL<4329> A_IWL<4328> A_IWL<4327> A_IWL<4326> A_IWL<4325> A_IWL<4324> A_IWL<4323> A_IWL<4322> A_IWL<4321> A_IWL<4320> A_IWL<4319> A_IWL<4318> A_IWL<4317> A_IWL<4316> A_IWL<4315> A_IWL<4314> A_IWL<4313> A_IWL<4312> A_IWL<4311> A_IWL<4310> A_IWL<4309> A_IWL<4308> A_IWL<4307> A_IWL<4306> A_IWL<4305> A_IWL<4304> A_IWL<4303> A_IWL<4302> A_IWL<4301> A_IWL<4300> A_IWL<4299> A_IWL<4298> A_IWL<4297> A_IWL<4296> A_IWL<4295> A_IWL<4294> A_IWL<4293> A_IWL<4292> A_IWL<4291> A_IWL<4290> A_IWL<4289> A_IWL<4288> A_IWL<4287> A_IWL<4286> A_IWL<4285> A_IWL<4284> A_IWL<4283> A_IWL<4282> A_IWL<4281> A_IWL<4280> A_IWL<4279> A_IWL<4278> A_IWL<4277> A_IWL<4276> A_IWL<4275> A_IWL<4274> A_IWL<4273> A_IWL<4272> A_IWL<4271> A_IWL<4270> A_IWL<4269> A_IWL<4268> A_IWL<4267> A_IWL<4266> A_IWL<4265> A_IWL<4264> A_IWL<4263> A_IWL<4262> A_IWL<4261> A_IWL<4260> A_IWL<4259> A_IWL<4258> A_IWL<4257> A_IWL<4256> A_IWL<4255> A_IWL<4254> A_IWL<4253> A_IWL<4252> A_IWL<4251> A_IWL<4250> A_IWL<4249> A_IWL<4248> A_IWL<4247> A_IWL<4246> A_IWL<4245> A_IWL<4244> A_IWL<4243> A_IWL<4242> A_IWL<4241> A_IWL<4240> A_IWL<4239> A_IWL<4238> A_IWL<4237> A_IWL<4236> A_IWL<4235> A_IWL<4234> A_IWL<4233> A_IWL<4232> A_IWL<4231> A_IWL<4230> A_IWL<4229> A_IWL<4228> A_IWL<4227> A_IWL<4226> A_IWL<4225> A_IWL<4224> A_IWL<4223> A_IWL<4222> A_IWL<4221> A_IWL<4220> A_IWL<4219> A_IWL<4218> A_IWL<4217> A_IWL<4216> A_IWL<4215> A_IWL<4214> A_IWL<4213> A_IWL<4212> A_IWL<4211> A_IWL<4210> A_IWL<4209> A_IWL<4208> A_IWL<4207> A_IWL<4206> A_IWL<4205> A_IWL<4204> A_IWL<4203> A_IWL<4202> A_IWL<4201> A_IWL<4200> A_IWL<4199> A_IWL<4198> A_IWL<4197> A_IWL<4196> A_IWL<4195> A_IWL<4194> A_IWL<4193> A_IWL<4192> A_IWL<4191> A_IWL<4190> A_IWL<4189> A_IWL<4188> A_IWL<4187> A_IWL<4186> A_IWL<4185> A_IWL<4184> A_IWL<4183> A_IWL<4182> A_IWL<4181> A_IWL<4180> A_IWL<4179> A_IWL<4178> A_IWL<4177> A_IWL<4176> A_IWL<4175> A_IWL<4174> A_IWL<4173> A_IWL<4172> A_IWL<4171> A_IWL<4170> A_IWL<4169> A_IWL<4168> A_IWL<4167> A_IWL<4166> A_IWL<4165> A_IWL<4164> A_IWL<4163> A_IWL<4162> A_IWL<4161> A_IWL<4160> A_IWL<4159> A_IWL<4158> A_IWL<4157> A_IWL<4156> A_IWL<4155> A_IWL<4154> A_IWL<4153> A_IWL<4152> A_IWL<4151> A_IWL<4150> A_IWL<4149> A_IWL<4148> A_IWL<4147> A_IWL<4146> A_IWL<4145> A_IWL<4144> A_IWL<4143> A_IWL<4142> A_IWL<4141> A_IWL<4140> A_IWL<4139> A_IWL<4138> A_IWL<4137> A_IWL<4136> A_IWL<4135> A_IWL<4134> A_IWL<4133> A_IWL<4132> A_IWL<4131> A_IWL<4130> A_IWL<4129> A_IWL<4128> A_IWL<4127> A_IWL<4126> A_IWL<4125> A_IWL<4124> A_IWL<4123> A_IWL<4122> A_IWL<4121> A_IWL<4120> A_IWL<4119> A_IWL<4118> A_IWL<4117> A_IWL<4116> A_IWL<4115> A_IWL<4114> A_IWL<4113> A_IWL<4112> A_IWL<4111> A_IWL<4110> A_IWL<4109> A_IWL<4108> A_IWL<4107> A_IWL<4106> A_IWL<4105> A_IWL<4104> A_IWL<4103> A_IWL<4102> A_IWL<4101> A_IWL<4100> A_IWL<4099> A_IWL<4098> A_IWL<4097> A_IWL<4096> A_IWL<4607> A_IWL<4606> A_IWL<4605> A_IWL<4604> A_IWL<4603> A_IWL<4602> A_IWL<4601> A_IWL<4600> A_IWL<4599> A_IWL<4598> A_IWL<4597> A_IWL<4596> A_IWL<4595> A_IWL<4594> A_IWL<4593> A_IWL<4592> A_IWL<4591> A_IWL<4590> A_IWL<4589> A_IWL<4588> A_IWL<4587> A_IWL<4586> A_IWL<4585> A_IWL<4584> A_IWL<4583> A_IWL<4582> A_IWL<4581> A_IWL<4580> A_IWL<4579> A_IWL<4578> A_IWL<4577> A_IWL<4576> A_IWL<4575> A_IWL<4574> A_IWL<4573> A_IWL<4572> A_IWL<4571> A_IWL<4570> A_IWL<4569> A_IWL<4568> A_IWL<4567> A_IWL<4566> A_IWL<4565> A_IWL<4564> A_IWL<4563> A_IWL<4562> A_IWL<4561> A_IWL<4560> A_IWL<4559> A_IWL<4558> A_IWL<4557> A_IWL<4556> A_IWL<4555> A_IWL<4554> A_IWL<4553> A_IWL<4552> A_IWL<4551> A_IWL<4550> A_IWL<4549> A_IWL<4548> A_IWL<4547> A_IWL<4546> A_IWL<4545> A_IWL<4544> A_IWL<4543> A_IWL<4542> A_IWL<4541> A_IWL<4540> A_IWL<4539> A_IWL<4538> A_IWL<4537> A_IWL<4536> A_IWL<4535> A_IWL<4534> A_IWL<4533> A_IWL<4532> A_IWL<4531> A_IWL<4530> A_IWL<4529> A_IWL<4528> A_IWL<4527> A_IWL<4526> A_IWL<4525> A_IWL<4524> A_IWL<4523> A_IWL<4522> A_IWL<4521> A_IWL<4520> A_IWL<4519> A_IWL<4518> A_IWL<4517> A_IWL<4516> A_IWL<4515> A_IWL<4514> A_IWL<4513> A_IWL<4512> A_IWL<4511> A_IWL<4510> A_IWL<4509> A_IWL<4508> A_IWL<4507> A_IWL<4506> A_IWL<4505> A_IWL<4504> A_IWL<4503> A_IWL<4502> A_IWL<4501> A_IWL<4500> A_IWL<4499> A_IWL<4498> A_IWL<4497> A_IWL<4496> A_IWL<4495> A_IWL<4494> A_IWL<4493> A_IWL<4492> A_IWL<4491> A_IWL<4490> A_IWL<4489> A_IWL<4488> A_IWL<4487> A_IWL<4486> A_IWL<4485> A_IWL<4484> A_IWL<4483> A_IWL<4482> A_IWL<4481> A_IWL<4480> A_IWL<4479> A_IWL<4478> A_IWL<4477> A_IWL<4476> A_IWL<4475> A_IWL<4474> A_IWL<4473> A_IWL<4472> A_IWL<4471> A_IWL<4470> A_IWL<4469> A_IWL<4468> A_IWL<4467> A_IWL<4466> A_IWL<4465> A_IWL<4464> A_IWL<4463> A_IWL<4462> A_IWL<4461> A_IWL<4460> A_IWL<4459> A_IWL<4458> A_IWL<4457> A_IWL<4456> A_IWL<4455> A_IWL<4454> A_IWL<4453> A_IWL<4452> A_IWL<4451> A_IWL<4450> A_IWL<4449> A_IWL<4448> A_IWL<4447> A_IWL<4446> A_IWL<4445> A_IWL<4444> A_IWL<4443> A_IWL<4442> A_IWL<4441> A_IWL<4440> A_IWL<4439> A_IWL<4438> A_IWL<4437> A_IWL<4436> A_IWL<4435> A_IWL<4434> A_IWL<4433> A_IWL<4432> A_IWL<4431> A_IWL<4430> A_IWL<4429> A_IWL<4428> A_IWL<4427> A_IWL<4426> A_IWL<4425> A_IWL<4424> A_IWL<4423> A_IWL<4422> A_IWL<4421> A_IWL<4420> A_IWL<4419> A_IWL<4418> A_IWL<4417> A_IWL<4416> A_IWL<4415> A_IWL<4414> A_IWL<4413> A_IWL<4412> A_IWL<4411> A_IWL<4410> A_IWL<4409> A_IWL<4408> A_IWL<4407> A_IWL<4406> A_IWL<4405> A_IWL<4404> A_IWL<4403> A_IWL<4402> A_IWL<4401> A_IWL<4400> A_IWL<4399> A_IWL<4398> A_IWL<4397> A_IWL<4396> A_IWL<4395> A_IWL<4394> A_IWL<4393> A_IWL<4392> A_IWL<4391> A_IWL<4390> A_IWL<4389> A_IWL<4388> A_IWL<4387> A_IWL<4386> A_IWL<4385> A_IWL<4384> A_IWL<4383> A_IWL<4382> A_IWL<4381> A_IWL<4380> A_IWL<4379> A_IWL<4378> A_IWL<4377> A_IWL<4376> A_IWL<4375> A_IWL<4374> A_IWL<4373> A_IWL<4372> A_IWL<4371> A_IWL<4370> A_IWL<4369> A_IWL<4368> A_IWL<4367> A_IWL<4366> A_IWL<4365> A_IWL<4364> A_IWL<4363> A_IWL<4362> A_IWL<4361> A_IWL<4360> A_IWL<4359> A_IWL<4358> A_IWL<4357> A_IWL<4356> A_IWL<4355> A_IWL<4354> A_IWL<4353> A_IWL<4352> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<16> A_BLC<33> A_BLC<32> A_BLC_TOP<33> A_BLC_TOP<32> A_BLT<33> A_BLT<32> A_BLT_TOP<33> A_BLT_TOP<32> A_IWL<4095> A_IWL<4094> A_IWL<4093> A_IWL<4092> A_IWL<4091> A_IWL<4090> A_IWL<4089> A_IWL<4088> A_IWL<4087> A_IWL<4086> A_IWL<4085> A_IWL<4084> A_IWL<4083> A_IWL<4082> A_IWL<4081> A_IWL<4080> A_IWL<4079> A_IWL<4078> A_IWL<4077> A_IWL<4076> A_IWL<4075> A_IWL<4074> A_IWL<4073> A_IWL<4072> A_IWL<4071> A_IWL<4070> A_IWL<4069> A_IWL<4068> A_IWL<4067> A_IWL<4066> A_IWL<4065> A_IWL<4064> A_IWL<4063> A_IWL<4062> A_IWL<4061> A_IWL<4060> A_IWL<4059> A_IWL<4058> A_IWL<4057> A_IWL<4056> A_IWL<4055> A_IWL<4054> A_IWL<4053> A_IWL<4052> A_IWL<4051> A_IWL<4050> A_IWL<4049> A_IWL<4048> A_IWL<4047> A_IWL<4046> A_IWL<4045> A_IWL<4044> A_IWL<4043> A_IWL<4042> A_IWL<4041> A_IWL<4040> A_IWL<4039> A_IWL<4038> A_IWL<4037> A_IWL<4036> A_IWL<4035> A_IWL<4034> A_IWL<4033> A_IWL<4032> A_IWL<4031> A_IWL<4030> A_IWL<4029> A_IWL<4028> A_IWL<4027> A_IWL<4026> A_IWL<4025> A_IWL<4024> A_IWL<4023> A_IWL<4022> A_IWL<4021> A_IWL<4020> A_IWL<4019> A_IWL<4018> A_IWL<4017> A_IWL<4016> A_IWL<4015> A_IWL<4014> A_IWL<4013> A_IWL<4012> A_IWL<4011> A_IWL<4010> A_IWL<4009> A_IWL<4008> A_IWL<4007> A_IWL<4006> A_IWL<4005> A_IWL<4004> A_IWL<4003> A_IWL<4002> A_IWL<4001> A_IWL<4000> A_IWL<3999> A_IWL<3998> A_IWL<3997> A_IWL<3996> A_IWL<3995> A_IWL<3994> A_IWL<3993> A_IWL<3992> A_IWL<3991> A_IWL<3990> A_IWL<3989> A_IWL<3988> A_IWL<3987> A_IWL<3986> A_IWL<3985> A_IWL<3984> A_IWL<3983> A_IWL<3982> A_IWL<3981> A_IWL<3980> A_IWL<3979> A_IWL<3978> A_IWL<3977> A_IWL<3976> A_IWL<3975> A_IWL<3974> A_IWL<3973> A_IWL<3972> A_IWL<3971> A_IWL<3970> A_IWL<3969> A_IWL<3968> A_IWL<3967> A_IWL<3966> A_IWL<3965> A_IWL<3964> A_IWL<3963> A_IWL<3962> A_IWL<3961> A_IWL<3960> A_IWL<3959> A_IWL<3958> A_IWL<3957> A_IWL<3956> A_IWL<3955> A_IWL<3954> A_IWL<3953> A_IWL<3952> A_IWL<3951> A_IWL<3950> A_IWL<3949> A_IWL<3948> A_IWL<3947> A_IWL<3946> A_IWL<3945> A_IWL<3944> A_IWL<3943> A_IWL<3942> A_IWL<3941> A_IWL<3940> A_IWL<3939> A_IWL<3938> A_IWL<3937> A_IWL<3936> A_IWL<3935> A_IWL<3934> A_IWL<3933> A_IWL<3932> A_IWL<3931> A_IWL<3930> A_IWL<3929> A_IWL<3928> A_IWL<3927> A_IWL<3926> A_IWL<3925> A_IWL<3924> A_IWL<3923> A_IWL<3922> A_IWL<3921> A_IWL<3920> A_IWL<3919> A_IWL<3918> A_IWL<3917> A_IWL<3916> A_IWL<3915> A_IWL<3914> A_IWL<3913> A_IWL<3912> A_IWL<3911> A_IWL<3910> A_IWL<3909> A_IWL<3908> A_IWL<3907> A_IWL<3906> A_IWL<3905> A_IWL<3904> A_IWL<3903> A_IWL<3902> A_IWL<3901> A_IWL<3900> A_IWL<3899> A_IWL<3898> A_IWL<3897> A_IWL<3896> A_IWL<3895> A_IWL<3894> A_IWL<3893> A_IWL<3892> A_IWL<3891> A_IWL<3890> A_IWL<3889> A_IWL<3888> A_IWL<3887> A_IWL<3886> A_IWL<3885> A_IWL<3884> A_IWL<3883> A_IWL<3882> A_IWL<3881> A_IWL<3880> A_IWL<3879> A_IWL<3878> A_IWL<3877> A_IWL<3876> A_IWL<3875> A_IWL<3874> A_IWL<3873> A_IWL<3872> A_IWL<3871> A_IWL<3870> A_IWL<3869> A_IWL<3868> A_IWL<3867> A_IWL<3866> A_IWL<3865> A_IWL<3864> A_IWL<3863> A_IWL<3862> A_IWL<3861> A_IWL<3860> A_IWL<3859> A_IWL<3858> A_IWL<3857> A_IWL<3856> A_IWL<3855> A_IWL<3854> A_IWL<3853> A_IWL<3852> A_IWL<3851> A_IWL<3850> A_IWL<3849> A_IWL<3848> A_IWL<3847> A_IWL<3846> A_IWL<3845> A_IWL<3844> A_IWL<3843> A_IWL<3842> A_IWL<3841> A_IWL<3840> A_IWL<4351> A_IWL<4350> A_IWL<4349> A_IWL<4348> A_IWL<4347> A_IWL<4346> A_IWL<4345> A_IWL<4344> A_IWL<4343> A_IWL<4342> A_IWL<4341> A_IWL<4340> A_IWL<4339> A_IWL<4338> A_IWL<4337> A_IWL<4336> A_IWL<4335> A_IWL<4334> A_IWL<4333> A_IWL<4332> A_IWL<4331> A_IWL<4330> A_IWL<4329> A_IWL<4328> A_IWL<4327> A_IWL<4326> A_IWL<4325> A_IWL<4324> A_IWL<4323> A_IWL<4322> A_IWL<4321> A_IWL<4320> A_IWL<4319> A_IWL<4318> A_IWL<4317> A_IWL<4316> A_IWL<4315> A_IWL<4314> A_IWL<4313> A_IWL<4312> A_IWL<4311> A_IWL<4310> A_IWL<4309> A_IWL<4308> A_IWL<4307> A_IWL<4306> A_IWL<4305> A_IWL<4304> A_IWL<4303> A_IWL<4302> A_IWL<4301> A_IWL<4300> A_IWL<4299> A_IWL<4298> A_IWL<4297> A_IWL<4296> A_IWL<4295> A_IWL<4294> A_IWL<4293> A_IWL<4292> A_IWL<4291> A_IWL<4290> A_IWL<4289> A_IWL<4288> A_IWL<4287> A_IWL<4286> A_IWL<4285> A_IWL<4284> A_IWL<4283> A_IWL<4282> A_IWL<4281> A_IWL<4280> A_IWL<4279> A_IWL<4278> A_IWL<4277> A_IWL<4276> A_IWL<4275> A_IWL<4274> A_IWL<4273> A_IWL<4272> A_IWL<4271> A_IWL<4270> A_IWL<4269> A_IWL<4268> A_IWL<4267> A_IWL<4266> A_IWL<4265> A_IWL<4264> A_IWL<4263> A_IWL<4262> A_IWL<4261> A_IWL<4260> A_IWL<4259> A_IWL<4258> A_IWL<4257> A_IWL<4256> A_IWL<4255> A_IWL<4254> A_IWL<4253> A_IWL<4252> A_IWL<4251> A_IWL<4250> A_IWL<4249> A_IWL<4248> A_IWL<4247> A_IWL<4246> A_IWL<4245> A_IWL<4244> A_IWL<4243> A_IWL<4242> A_IWL<4241> A_IWL<4240> A_IWL<4239> A_IWL<4238> A_IWL<4237> A_IWL<4236> A_IWL<4235> A_IWL<4234> A_IWL<4233> A_IWL<4232> A_IWL<4231> A_IWL<4230> A_IWL<4229> A_IWL<4228> A_IWL<4227> A_IWL<4226> A_IWL<4225> A_IWL<4224> A_IWL<4223> A_IWL<4222> A_IWL<4221> A_IWL<4220> A_IWL<4219> A_IWL<4218> A_IWL<4217> A_IWL<4216> A_IWL<4215> A_IWL<4214> A_IWL<4213> A_IWL<4212> A_IWL<4211> A_IWL<4210> A_IWL<4209> A_IWL<4208> A_IWL<4207> A_IWL<4206> A_IWL<4205> A_IWL<4204> A_IWL<4203> A_IWL<4202> A_IWL<4201> A_IWL<4200> A_IWL<4199> A_IWL<4198> A_IWL<4197> A_IWL<4196> A_IWL<4195> A_IWL<4194> A_IWL<4193> A_IWL<4192> A_IWL<4191> A_IWL<4190> A_IWL<4189> A_IWL<4188> A_IWL<4187> A_IWL<4186> A_IWL<4185> A_IWL<4184> A_IWL<4183> A_IWL<4182> A_IWL<4181> A_IWL<4180> A_IWL<4179> A_IWL<4178> A_IWL<4177> A_IWL<4176> A_IWL<4175> A_IWL<4174> A_IWL<4173> A_IWL<4172> A_IWL<4171> A_IWL<4170> A_IWL<4169> A_IWL<4168> A_IWL<4167> A_IWL<4166> A_IWL<4165> A_IWL<4164> A_IWL<4163> A_IWL<4162> A_IWL<4161> A_IWL<4160> A_IWL<4159> A_IWL<4158> A_IWL<4157> A_IWL<4156> A_IWL<4155> A_IWL<4154> A_IWL<4153> A_IWL<4152> A_IWL<4151> A_IWL<4150> A_IWL<4149> A_IWL<4148> A_IWL<4147> A_IWL<4146> A_IWL<4145> A_IWL<4144> A_IWL<4143> A_IWL<4142> A_IWL<4141> A_IWL<4140> A_IWL<4139> A_IWL<4138> A_IWL<4137> A_IWL<4136> A_IWL<4135> A_IWL<4134> A_IWL<4133> A_IWL<4132> A_IWL<4131> A_IWL<4130> A_IWL<4129> A_IWL<4128> A_IWL<4127> A_IWL<4126> A_IWL<4125> A_IWL<4124> A_IWL<4123> A_IWL<4122> A_IWL<4121> A_IWL<4120> A_IWL<4119> A_IWL<4118> A_IWL<4117> A_IWL<4116> A_IWL<4115> A_IWL<4114> A_IWL<4113> A_IWL<4112> A_IWL<4111> A_IWL<4110> A_IWL<4109> A_IWL<4108> A_IWL<4107> A_IWL<4106> A_IWL<4105> A_IWL<4104> A_IWL<4103> A_IWL<4102> A_IWL<4101> A_IWL<4100> A_IWL<4099> A_IWL<4098> A_IWL<4097> A_IWL<4096> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<15> A_BLC<31> A_BLC<30> A_BLC_TOP<31> A_BLC_TOP<30> A_BLT<31> A_BLT<30> A_BLT_TOP<31> A_BLT_TOP<30> A_IWL<3839> A_IWL<3838> A_IWL<3837> A_IWL<3836> A_IWL<3835> A_IWL<3834> A_IWL<3833> A_IWL<3832> A_IWL<3831> A_IWL<3830> A_IWL<3829> A_IWL<3828> A_IWL<3827> A_IWL<3826> A_IWL<3825> A_IWL<3824> A_IWL<3823> A_IWL<3822> A_IWL<3821> A_IWL<3820> A_IWL<3819> A_IWL<3818> A_IWL<3817> A_IWL<3816> A_IWL<3815> A_IWL<3814> A_IWL<3813> A_IWL<3812> A_IWL<3811> A_IWL<3810> A_IWL<3809> A_IWL<3808> A_IWL<3807> A_IWL<3806> A_IWL<3805> A_IWL<3804> A_IWL<3803> A_IWL<3802> A_IWL<3801> A_IWL<3800> A_IWL<3799> A_IWL<3798> A_IWL<3797> A_IWL<3796> A_IWL<3795> A_IWL<3794> A_IWL<3793> A_IWL<3792> A_IWL<3791> A_IWL<3790> A_IWL<3789> A_IWL<3788> A_IWL<3787> A_IWL<3786> A_IWL<3785> A_IWL<3784> A_IWL<3783> A_IWL<3782> A_IWL<3781> A_IWL<3780> A_IWL<3779> A_IWL<3778> A_IWL<3777> A_IWL<3776> A_IWL<3775> A_IWL<3774> A_IWL<3773> A_IWL<3772> A_IWL<3771> A_IWL<3770> A_IWL<3769> A_IWL<3768> A_IWL<3767> A_IWL<3766> A_IWL<3765> A_IWL<3764> A_IWL<3763> A_IWL<3762> A_IWL<3761> A_IWL<3760> A_IWL<3759> A_IWL<3758> A_IWL<3757> A_IWL<3756> A_IWL<3755> A_IWL<3754> A_IWL<3753> A_IWL<3752> A_IWL<3751> A_IWL<3750> A_IWL<3749> A_IWL<3748> A_IWL<3747> A_IWL<3746> A_IWL<3745> A_IWL<3744> A_IWL<3743> A_IWL<3742> A_IWL<3741> A_IWL<3740> A_IWL<3739> A_IWL<3738> A_IWL<3737> A_IWL<3736> A_IWL<3735> A_IWL<3734> A_IWL<3733> A_IWL<3732> A_IWL<3731> A_IWL<3730> A_IWL<3729> A_IWL<3728> A_IWL<3727> A_IWL<3726> A_IWL<3725> A_IWL<3724> A_IWL<3723> A_IWL<3722> A_IWL<3721> A_IWL<3720> A_IWL<3719> A_IWL<3718> A_IWL<3717> A_IWL<3716> A_IWL<3715> A_IWL<3714> A_IWL<3713> A_IWL<3712> A_IWL<3711> A_IWL<3710> A_IWL<3709> A_IWL<3708> A_IWL<3707> A_IWL<3706> A_IWL<3705> A_IWL<3704> A_IWL<3703> A_IWL<3702> A_IWL<3701> A_IWL<3700> A_IWL<3699> A_IWL<3698> A_IWL<3697> A_IWL<3696> A_IWL<3695> A_IWL<3694> A_IWL<3693> A_IWL<3692> A_IWL<3691> A_IWL<3690> A_IWL<3689> A_IWL<3688> A_IWL<3687> A_IWL<3686> A_IWL<3685> A_IWL<3684> A_IWL<3683> A_IWL<3682> A_IWL<3681> A_IWL<3680> A_IWL<3679> A_IWL<3678> A_IWL<3677> A_IWL<3676> A_IWL<3675> A_IWL<3674> A_IWL<3673> A_IWL<3672> A_IWL<3671> A_IWL<3670> A_IWL<3669> A_IWL<3668> A_IWL<3667> A_IWL<3666> A_IWL<3665> A_IWL<3664> A_IWL<3663> A_IWL<3662> A_IWL<3661> A_IWL<3660> A_IWL<3659> A_IWL<3658> A_IWL<3657> A_IWL<3656> A_IWL<3655> A_IWL<3654> A_IWL<3653> A_IWL<3652> A_IWL<3651> A_IWL<3650> A_IWL<3649> A_IWL<3648> A_IWL<3647> A_IWL<3646> A_IWL<3645> A_IWL<3644> A_IWL<3643> A_IWL<3642> A_IWL<3641> A_IWL<3640> A_IWL<3639> A_IWL<3638> A_IWL<3637> A_IWL<3636> A_IWL<3635> A_IWL<3634> A_IWL<3633> A_IWL<3632> A_IWL<3631> A_IWL<3630> A_IWL<3629> A_IWL<3628> A_IWL<3627> A_IWL<3626> A_IWL<3625> A_IWL<3624> A_IWL<3623> A_IWL<3622> A_IWL<3621> A_IWL<3620> A_IWL<3619> A_IWL<3618> A_IWL<3617> A_IWL<3616> A_IWL<3615> A_IWL<3614> A_IWL<3613> A_IWL<3612> A_IWL<3611> A_IWL<3610> A_IWL<3609> A_IWL<3608> A_IWL<3607> A_IWL<3606> A_IWL<3605> A_IWL<3604> A_IWL<3603> A_IWL<3602> A_IWL<3601> A_IWL<3600> A_IWL<3599> A_IWL<3598> A_IWL<3597> A_IWL<3596> A_IWL<3595> A_IWL<3594> A_IWL<3593> A_IWL<3592> A_IWL<3591> A_IWL<3590> A_IWL<3589> A_IWL<3588> A_IWL<3587> A_IWL<3586> A_IWL<3585> A_IWL<3584> A_IWL<4095> A_IWL<4094> A_IWL<4093> A_IWL<4092> A_IWL<4091> A_IWL<4090> A_IWL<4089> A_IWL<4088> A_IWL<4087> A_IWL<4086> A_IWL<4085> A_IWL<4084> A_IWL<4083> A_IWL<4082> A_IWL<4081> A_IWL<4080> A_IWL<4079> A_IWL<4078> A_IWL<4077> A_IWL<4076> A_IWL<4075> A_IWL<4074> A_IWL<4073> A_IWL<4072> A_IWL<4071> A_IWL<4070> A_IWL<4069> A_IWL<4068> A_IWL<4067> A_IWL<4066> A_IWL<4065> A_IWL<4064> A_IWL<4063> A_IWL<4062> A_IWL<4061> A_IWL<4060> A_IWL<4059> A_IWL<4058> A_IWL<4057> A_IWL<4056> A_IWL<4055> A_IWL<4054> A_IWL<4053> A_IWL<4052> A_IWL<4051> A_IWL<4050> A_IWL<4049> A_IWL<4048> A_IWL<4047> A_IWL<4046> A_IWL<4045> A_IWL<4044> A_IWL<4043> A_IWL<4042> A_IWL<4041> A_IWL<4040> A_IWL<4039> A_IWL<4038> A_IWL<4037> A_IWL<4036> A_IWL<4035> A_IWL<4034> A_IWL<4033> A_IWL<4032> A_IWL<4031> A_IWL<4030> A_IWL<4029> A_IWL<4028> A_IWL<4027> A_IWL<4026> A_IWL<4025> A_IWL<4024> A_IWL<4023> A_IWL<4022> A_IWL<4021> A_IWL<4020> A_IWL<4019> A_IWL<4018> A_IWL<4017> A_IWL<4016> A_IWL<4015> A_IWL<4014> A_IWL<4013> A_IWL<4012> A_IWL<4011> A_IWL<4010> A_IWL<4009> A_IWL<4008> A_IWL<4007> A_IWL<4006> A_IWL<4005> A_IWL<4004> A_IWL<4003> A_IWL<4002> A_IWL<4001> A_IWL<4000> A_IWL<3999> A_IWL<3998> A_IWL<3997> A_IWL<3996> A_IWL<3995> A_IWL<3994> A_IWL<3993> A_IWL<3992> A_IWL<3991> A_IWL<3990> A_IWL<3989> A_IWL<3988> A_IWL<3987> A_IWL<3986> A_IWL<3985> A_IWL<3984> A_IWL<3983> A_IWL<3982> A_IWL<3981> A_IWL<3980> A_IWL<3979> A_IWL<3978> A_IWL<3977> A_IWL<3976> A_IWL<3975> A_IWL<3974> A_IWL<3973> A_IWL<3972> A_IWL<3971> A_IWL<3970> A_IWL<3969> A_IWL<3968> A_IWL<3967> A_IWL<3966> A_IWL<3965> A_IWL<3964> A_IWL<3963> A_IWL<3962> A_IWL<3961> A_IWL<3960> A_IWL<3959> A_IWL<3958> A_IWL<3957> A_IWL<3956> A_IWL<3955> A_IWL<3954> A_IWL<3953> A_IWL<3952> A_IWL<3951> A_IWL<3950> A_IWL<3949> A_IWL<3948> A_IWL<3947> A_IWL<3946> A_IWL<3945> A_IWL<3944> A_IWL<3943> A_IWL<3942> A_IWL<3941> A_IWL<3940> A_IWL<3939> A_IWL<3938> A_IWL<3937> A_IWL<3936> A_IWL<3935> A_IWL<3934> A_IWL<3933> A_IWL<3932> A_IWL<3931> A_IWL<3930> A_IWL<3929> A_IWL<3928> A_IWL<3927> A_IWL<3926> A_IWL<3925> A_IWL<3924> A_IWL<3923> A_IWL<3922> A_IWL<3921> A_IWL<3920> A_IWL<3919> A_IWL<3918> A_IWL<3917> A_IWL<3916> A_IWL<3915> A_IWL<3914> A_IWL<3913> A_IWL<3912> A_IWL<3911> A_IWL<3910> A_IWL<3909> A_IWL<3908> A_IWL<3907> A_IWL<3906> A_IWL<3905> A_IWL<3904> A_IWL<3903> A_IWL<3902> A_IWL<3901> A_IWL<3900> A_IWL<3899> A_IWL<3898> A_IWL<3897> A_IWL<3896> A_IWL<3895> A_IWL<3894> A_IWL<3893> A_IWL<3892> A_IWL<3891> A_IWL<3890> A_IWL<3889> A_IWL<3888> A_IWL<3887> A_IWL<3886> A_IWL<3885> A_IWL<3884> A_IWL<3883> A_IWL<3882> A_IWL<3881> A_IWL<3880> A_IWL<3879> A_IWL<3878> A_IWL<3877> A_IWL<3876> A_IWL<3875> A_IWL<3874> A_IWL<3873> A_IWL<3872> A_IWL<3871> A_IWL<3870> A_IWL<3869> A_IWL<3868> A_IWL<3867> A_IWL<3866> A_IWL<3865> A_IWL<3864> A_IWL<3863> A_IWL<3862> A_IWL<3861> A_IWL<3860> A_IWL<3859> A_IWL<3858> A_IWL<3857> A_IWL<3856> A_IWL<3855> A_IWL<3854> A_IWL<3853> A_IWL<3852> A_IWL<3851> A_IWL<3850> A_IWL<3849> A_IWL<3848> A_IWL<3847> A_IWL<3846> A_IWL<3845> A_IWL<3844> A_IWL<3843> A_IWL<3842> A_IWL<3841> A_IWL<3840> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<14> A_BLC<29> A_BLC<28> A_BLC_TOP<29> A_BLC_TOP<28> A_BLT<29> A_BLT<28> A_BLT_TOP<29> A_BLT_TOP<28> A_IWL<3583> A_IWL<3582> A_IWL<3581> A_IWL<3580> A_IWL<3579> A_IWL<3578> A_IWL<3577> A_IWL<3576> A_IWL<3575> A_IWL<3574> A_IWL<3573> A_IWL<3572> A_IWL<3571> A_IWL<3570> A_IWL<3569> A_IWL<3568> A_IWL<3567> A_IWL<3566> A_IWL<3565> A_IWL<3564> A_IWL<3563> A_IWL<3562> A_IWL<3561> A_IWL<3560> A_IWL<3559> A_IWL<3558> A_IWL<3557> A_IWL<3556> A_IWL<3555> A_IWL<3554> A_IWL<3553> A_IWL<3552> A_IWL<3551> A_IWL<3550> A_IWL<3549> A_IWL<3548> A_IWL<3547> A_IWL<3546> A_IWL<3545> A_IWL<3544> A_IWL<3543> A_IWL<3542> A_IWL<3541> A_IWL<3540> A_IWL<3539> A_IWL<3538> A_IWL<3537> A_IWL<3536> A_IWL<3535> A_IWL<3534> A_IWL<3533> A_IWL<3532> A_IWL<3531> A_IWL<3530> A_IWL<3529> A_IWL<3528> A_IWL<3527> A_IWL<3526> A_IWL<3525> A_IWL<3524> A_IWL<3523> A_IWL<3522> A_IWL<3521> A_IWL<3520> A_IWL<3519> A_IWL<3518> A_IWL<3517> A_IWL<3516> A_IWL<3515> A_IWL<3514> A_IWL<3513> A_IWL<3512> A_IWL<3511> A_IWL<3510> A_IWL<3509> A_IWL<3508> A_IWL<3507> A_IWL<3506> A_IWL<3505> A_IWL<3504> A_IWL<3503> A_IWL<3502> A_IWL<3501> A_IWL<3500> A_IWL<3499> A_IWL<3498> A_IWL<3497> A_IWL<3496> A_IWL<3495> A_IWL<3494> A_IWL<3493> A_IWL<3492> A_IWL<3491> A_IWL<3490> A_IWL<3489> A_IWL<3488> A_IWL<3487> A_IWL<3486> A_IWL<3485> A_IWL<3484> A_IWL<3483> A_IWL<3482> A_IWL<3481> A_IWL<3480> A_IWL<3479> A_IWL<3478> A_IWL<3477> A_IWL<3476> A_IWL<3475> A_IWL<3474> A_IWL<3473> A_IWL<3472> A_IWL<3471> A_IWL<3470> A_IWL<3469> A_IWL<3468> A_IWL<3467> A_IWL<3466> A_IWL<3465> A_IWL<3464> A_IWL<3463> A_IWL<3462> A_IWL<3461> A_IWL<3460> A_IWL<3459> A_IWL<3458> A_IWL<3457> A_IWL<3456> A_IWL<3455> A_IWL<3454> A_IWL<3453> A_IWL<3452> A_IWL<3451> A_IWL<3450> A_IWL<3449> A_IWL<3448> A_IWL<3447> A_IWL<3446> A_IWL<3445> A_IWL<3444> A_IWL<3443> A_IWL<3442> A_IWL<3441> A_IWL<3440> A_IWL<3439> A_IWL<3438> A_IWL<3437> A_IWL<3436> A_IWL<3435> A_IWL<3434> A_IWL<3433> A_IWL<3432> A_IWL<3431> A_IWL<3430> A_IWL<3429> A_IWL<3428> A_IWL<3427> A_IWL<3426> A_IWL<3425> A_IWL<3424> A_IWL<3423> A_IWL<3422> A_IWL<3421> A_IWL<3420> A_IWL<3419> A_IWL<3418> A_IWL<3417> A_IWL<3416> A_IWL<3415> A_IWL<3414> A_IWL<3413> A_IWL<3412> A_IWL<3411> A_IWL<3410> A_IWL<3409> A_IWL<3408> A_IWL<3407> A_IWL<3406> A_IWL<3405> A_IWL<3404> A_IWL<3403> A_IWL<3402> A_IWL<3401> A_IWL<3400> A_IWL<3399> A_IWL<3398> A_IWL<3397> A_IWL<3396> A_IWL<3395> A_IWL<3394> A_IWL<3393> A_IWL<3392> A_IWL<3391> A_IWL<3390> A_IWL<3389> A_IWL<3388> A_IWL<3387> A_IWL<3386> A_IWL<3385> A_IWL<3384> A_IWL<3383> A_IWL<3382> A_IWL<3381> A_IWL<3380> A_IWL<3379> A_IWL<3378> A_IWL<3377> A_IWL<3376> A_IWL<3375> A_IWL<3374> A_IWL<3373> A_IWL<3372> A_IWL<3371> A_IWL<3370> A_IWL<3369> A_IWL<3368> A_IWL<3367> A_IWL<3366> A_IWL<3365> A_IWL<3364> A_IWL<3363> A_IWL<3362> A_IWL<3361> A_IWL<3360> A_IWL<3359> A_IWL<3358> A_IWL<3357> A_IWL<3356> A_IWL<3355> A_IWL<3354> A_IWL<3353> A_IWL<3352> A_IWL<3351> A_IWL<3350> A_IWL<3349> A_IWL<3348> A_IWL<3347> A_IWL<3346> A_IWL<3345> A_IWL<3344> A_IWL<3343> A_IWL<3342> A_IWL<3341> A_IWL<3340> A_IWL<3339> A_IWL<3338> A_IWL<3337> A_IWL<3336> A_IWL<3335> A_IWL<3334> A_IWL<3333> A_IWL<3332> A_IWL<3331> A_IWL<3330> A_IWL<3329> A_IWL<3328> A_IWL<3839> A_IWL<3838> A_IWL<3837> A_IWL<3836> A_IWL<3835> A_IWL<3834> A_IWL<3833> A_IWL<3832> A_IWL<3831> A_IWL<3830> A_IWL<3829> A_IWL<3828> A_IWL<3827> A_IWL<3826> A_IWL<3825> A_IWL<3824> A_IWL<3823> A_IWL<3822> A_IWL<3821> A_IWL<3820> A_IWL<3819> A_IWL<3818> A_IWL<3817> A_IWL<3816> A_IWL<3815> A_IWL<3814> A_IWL<3813> A_IWL<3812> A_IWL<3811> A_IWL<3810> A_IWL<3809> A_IWL<3808> A_IWL<3807> A_IWL<3806> A_IWL<3805> A_IWL<3804> A_IWL<3803> A_IWL<3802> A_IWL<3801> A_IWL<3800> A_IWL<3799> A_IWL<3798> A_IWL<3797> A_IWL<3796> A_IWL<3795> A_IWL<3794> A_IWL<3793> A_IWL<3792> A_IWL<3791> A_IWL<3790> A_IWL<3789> A_IWL<3788> A_IWL<3787> A_IWL<3786> A_IWL<3785> A_IWL<3784> A_IWL<3783> A_IWL<3782> A_IWL<3781> A_IWL<3780> A_IWL<3779> A_IWL<3778> A_IWL<3777> A_IWL<3776> A_IWL<3775> A_IWL<3774> A_IWL<3773> A_IWL<3772> A_IWL<3771> A_IWL<3770> A_IWL<3769> A_IWL<3768> A_IWL<3767> A_IWL<3766> A_IWL<3765> A_IWL<3764> A_IWL<3763> A_IWL<3762> A_IWL<3761> A_IWL<3760> A_IWL<3759> A_IWL<3758> A_IWL<3757> A_IWL<3756> A_IWL<3755> A_IWL<3754> A_IWL<3753> A_IWL<3752> A_IWL<3751> A_IWL<3750> A_IWL<3749> A_IWL<3748> A_IWL<3747> A_IWL<3746> A_IWL<3745> A_IWL<3744> A_IWL<3743> A_IWL<3742> A_IWL<3741> A_IWL<3740> A_IWL<3739> A_IWL<3738> A_IWL<3737> A_IWL<3736> A_IWL<3735> A_IWL<3734> A_IWL<3733> A_IWL<3732> A_IWL<3731> A_IWL<3730> A_IWL<3729> A_IWL<3728> A_IWL<3727> A_IWL<3726> A_IWL<3725> A_IWL<3724> A_IWL<3723> A_IWL<3722> A_IWL<3721> A_IWL<3720> A_IWL<3719> A_IWL<3718> A_IWL<3717> A_IWL<3716> A_IWL<3715> A_IWL<3714> A_IWL<3713> A_IWL<3712> A_IWL<3711> A_IWL<3710> A_IWL<3709> A_IWL<3708> A_IWL<3707> A_IWL<3706> A_IWL<3705> A_IWL<3704> A_IWL<3703> A_IWL<3702> A_IWL<3701> A_IWL<3700> A_IWL<3699> A_IWL<3698> A_IWL<3697> A_IWL<3696> A_IWL<3695> A_IWL<3694> A_IWL<3693> A_IWL<3692> A_IWL<3691> A_IWL<3690> A_IWL<3689> A_IWL<3688> A_IWL<3687> A_IWL<3686> A_IWL<3685> A_IWL<3684> A_IWL<3683> A_IWL<3682> A_IWL<3681> A_IWL<3680> A_IWL<3679> A_IWL<3678> A_IWL<3677> A_IWL<3676> A_IWL<3675> A_IWL<3674> A_IWL<3673> A_IWL<3672> A_IWL<3671> A_IWL<3670> A_IWL<3669> A_IWL<3668> A_IWL<3667> A_IWL<3666> A_IWL<3665> A_IWL<3664> A_IWL<3663> A_IWL<3662> A_IWL<3661> A_IWL<3660> A_IWL<3659> A_IWL<3658> A_IWL<3657> A_IWL<3656> A_IWL<3655> A_IWL<3654> A_IWL<3653> A_IWL<3652> A_IWL<3651> A_IWL<3650> A_IWL<3649> A_IWL<3648> A_IWL<3647> A_IWL<3646> A_IWL<3645> A_IWL<3644> A_IWL<3643> A_IWL<3642> A_IWL<3641> A_IWL<3640> A_IWL<3639> A_IWL<3638> A_IWL<3637> A_IWL<3636> A_IWL<3635> A_IWL<3634> A_IWL<3633> A_IWL<3632> A_IWL<3631> A_IWL<3630> A_IWL<3629> A_IWL<3628> A_IWL<3627> A_IWL<3626> A_IWL<3625> A_IWL<3624> A_IWL<3623> A_IWL<3622> A_IWL<3621> A_IWL<3620> A_IWL<3619> A_IWL<3618> A_IWL<3617> A_IWL<3616> A_IWL<3615> A_IWL<3614> A_IWL<3613> A_IWL<3612> A_IWL<3611> A_IWL<3610> A_IWL<3609> A_IWL<3608> A_IWL<3607> A_IWL<3606> A_IWL<3605> A_IWL<3604> A_IWL<3603> A_IWL<3602> A_IWL<3601> A_IWL<3600> A_IWL<3599> A_IWL<3598> A_IWL<3597> A_IWL<3596> A_IWL<3595> A_IWL<3594> A_IWL<3593> A_IWL<3592> A_IWL<3591> A_IWL<3590> A_IWL<3589> A_IWL<3588> A_IWL<3587> A_IWL<3586> A_IWL<3585> A_IWL<3584> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<13> A_BLC<27> A_BLC<26> A_BLC_TOP<27> A_BLC_TOP<26> A_BLT<27> A_BLT<26> A_BLT_TOP<27> A_BLT_TOP<26> A_IWL<3327> A_IWL<3326> A_IWL<3325> A_IWL<3324> A_IWL<3323> A_IWL<3322> A_IWL<3321> A_IWL<3320> A_IWL<3319> A_IWL<3318> A_IWL<3317> A_IWL<3316> A_IWL<3315> A_IWL<3314> A_IWL<3313> A_IWL<3312> A_IWL<3311> A_IWL<3310> A_IWL<3309> A_IWL<3308> A_IWL<3307> A_IWL<3306> A_IWL<3305> A_IWL<3304> A_IWL<3303> A_IWL<3302> A_IWL<3301> A_IWL<3300> A_IWL<3299> A_IWL<3298> A_IWL<3297> A_IWL<3296> A_IWL<3295> A_IWL<3294> A_IWL<3293> A_IWL<3292> A_IWL<3291> A_IWL<3290> A_IWL<3289> A_IWL<3288> A_IWL<3287> A_IWL<3286> A_IWL<3285> A_IWL<3284> A_IWL<3283> A_IWL<3282> A_IWL<3281> A_IWL<3280> A_IWL<3279> A_IWL<3278> A_IWL<3277> A_IWL<3276> A_IWL<3275> A_IWL<3274> A_IWL<3273> A_IWL<3272> A_IWL<3271> A_IWL<3270> A_IWL<3269> A_IWL<3268> A_IWL<3267> A_IWL<3266> A_IWL<3265> A_IWL<3264> A_IWL<3263> A_IWL<3262> A_IWL<3261> A_IWL<3260> A_IWL<3259> A_IWL<3258> A_IWL<3257> A_IWL<3256> A_IWL<3255> A_IWL<3254> A_IWL<3253> A_IWL<3252> A_IWL<3251> A_IWL<3250> A_IWL<3249> A_IWL<3248> A_IWL<3247> A_IWL<3246> A_IWL<3245> A_IWL<3244> A_IWL<3243> A_IWL<3242> A_IWL<3241> A_IWL<3240> A_IWL<3239> A_IWL<3238> A_IWL<3237> A_IWL<3236> A_IWL<3235> A_IWL<3234> A_IWL<3233> A_IWL<3232> A_IWL<3231> A_IWL<3230> A_IWL<3229> A_IWL<3228> A_IWL<3227> A_IWL<3226> A_IWL<3225> A_IWL<3224> A_IWL<3223> A_IWL<3222> A_IWL<3221> A_IWL<3220> A_IWL<3219> A_IWL<3218> A_IWL<3217> A_IWL<3216> A_IWL<3215> A_IWL<3214> A_IWL<3213> A_IWL<3212> A_IWL<3211> A_IWL<3210> A_IWL<3209> A_IWL<3208> A_IWL<3207> A_IWL<3206> A_IWL<3205> A_IWL<3204> A_IWL<3203> A_IWL<3202> A_IWL<3201> A_IWL<3200> A_IWL<3199> A_IWL<3198> A_IWL<3197> A_IWL<3196> A_IWL<3195> A_IWL<3194> A_IWL<3193> A_IWL<3192> A_IWL<3191> A_IWL<3190> A_IWL<3189> A_IWL<3188> A_IWL<3187> A_IWL<3186> A_IWL<3185> A_IWL<3184> A_IWL<3183> A_IWL<3182> A_IWL<3181> A_IWL<3180> A_IWL<3179> A_IWL<3178> A_IWL<3177> A_IWL<3176> A_IWL<3175> A_IWL<3174> A_IWL<3173> A_IWL<3172> A_IWL<3171> A_IWL<3170> A_IWL<3169> A_IWL<3168> A_IWL<3167> A_IWL<3166> A_IWL<3165> A_IWL<3164> A_IWL<3163> A_IWL<3162> A_IWL<3161> A_IWL<3160> A_IWL<3159> A_IWL<3158> A_IWL<3157> A_IWL<3156> A_IWL<3155> A_IWL<3154> A_IWL<3153> A_IWL<3152> A_IWL<3151> A_IWL<3150> A_IWL<3149> A_IWL<3148> A_IWL<3147> A_IWL<3146> A_IWL<3145> A_IWL<3144> A_IWL<3143> A_IWL<3142> A_IWL<3141> A_IWL<3140> A_IWL<3139> A_IWL<3138> A_IWL<3137> A_IWL<3136> A_IWL<3135> A_IWL<3134> A_IWL<3133> A_IWL<3132> A_IWL<3131> A_IWL<3130> A_IWL<3129> A_IWL<3128> A_IWL<3127> A_IWL<3126> A_IWL<3125> A_IWL<3124> A_IWL<3123> A_IWL<3122> A_IWL<3121> A_IWL<3120> A_IWL<3119> A_IWL<3118> A_IWL<3117> A_IWL<3116> A_IWL<3115> A_IWL<3114> A_IWL<3113> A_IWL<3112> A_IWL<3111> A_IWL<3110> A_IWL<3109> A_IWL<3108> A_IWL<3107> A_IWL<3106> A_IWL<3105> A_IWL<3104> A_IWL<3103> A_IWL<3102> A_IWL<3101> A_IWL<3100> A_IWL<3099> A_IWL<3098> A_IWL<3097> A_IWL<3096> A_IWL<3095> A_IWL<3094> A_IWL<3093> A_IWL<3092> A_IWL<3091> A_IWL<3090> A_IWL<3089> A_IWL<3088> A_IWL<3087> A_IWL<3086> A_IWL<3085> A_IWL<3084> A_IWL<3083> A_IWL<3082> A_IWL<3081> A_IWL<3080> A_IWL<3079> A_IWL<3078> A_IWL<3077> A_IWL<3076> A_IWL<3075> A_IWL<3074> A_IWL<3073> A_IWL<3072> A_IWL<3583> A_IWL<3582> A_IWL<3581> A_IWL<3580> A_IWL<3579> A_IWL<3578> A_IWL<3577> A_IWL<3576> A_IWL<3575> A_IWL<3574> A_IWL<3573> A_IWL<3572> A_IWL<3571> A_IWL<3570> A_IWL<3569> A_IWL<3568> A_IWL<3567> A_IWL<3566> A_IWL<3565> A_IWL<3564> A_IWL<3563> A_IWL<3562> A_IWL<3561> A_IWL<3560> A_IWL<3559> A_IWL<3558> A_IWL<3557> A_IWL<3556> A_IWL<3555> A_IWL<3554> A_IWL<3553> A_IWL<3552> A_IWL<3551> A_IWL<3550> A_IWL<3549> A_IWL<3548> A_IWL<3547> A_IWL<3546> A_IWL<3545> A_IWL<3544> A_IWL<3543> A_IWL<3542> A_IWL<3541> A_IWL<3540> A_IWL<3539> A_IWL<3538> A_IWL<3537> A_IWL<3536> A_IWL<3535> A_IWL<3534> A_IWL<3533> A_IWL<3532> A_IWL<3531> A_IWL<3530> A_IWL<3529> A_IWL<3528> A_IWL<3527> A_IWL<3526> A_IWL<3525> A_IWL<3524> A_IWL<3523> A_IWL<3522> A_IWL<3521> A_IWL<3520> A_IWL<3519> A_IWL<3518> A_IWL<3517> A_IWL<3516> A_IWL<3515> A_IWL<3514> A_IWL<3513> A_IWL<3512> A_IWL<3511> A_IWL<3510> A_IWL<3509> A_IWL<3508> A_IWL<3507> A_IWL<3506> A_IWL<3505> A_IWL<3504> A_IWL<3503> A_IWL<3502> A_IWL<3501> A_IWL<3500> A_IWL<3499> A_IWL<3498> A_IWL<3497> A_IWL<3496> A_IWL<3495> A_IWL<3494> A_IWL<3493> A_IWL<3492> A_IWL<3491> A_IWL<3490> A_IWL<3489> A_IWL<3488> A_IWL<3487> A_IWL<3486> A_IWL<3485> A_IWL<3484> A_IWL<3483> A_IWL<3482> A_IWL<3481> A_IWL<3480> A_IWL<3479> A_IWL<3478> A_IWL<3477> A_IWL<3476> A_IWL<3475> A_IWL<3474> A_IWL<3473> A_IWL<3472> A_IWL<3471> A_IWL<3470> A_IWL<3469> A_IWL<3468> A_IWL<3467> A_IWL<3466> A_IWL<3465> A_IWL<3464> A_IWL<3463> A_IWL<3462> A_IWL<3461> A_IWL<3460> A_IWL<3459> A_IWL<3458> A_IWL<3457> A_IWL<3456> A_IWL<3455> A_IWL<3454> A_IWL<3453> A_IWL<3452> A_IWL<3451> A_IWL<3450> A_IWL<3449> A_IWL<3448> A_IWL<3447> A_IWL<3446> A_IWL<3445> A_IWL<3444> A_IWL<3443> A_IWL<3442> A_IWL<3441> A_IWL<3440> A_IWL<3439> A_IWL<3438> A_IWL<3437> A_IWL<3436> A_IWL<3435> A_IWL<3434> A_IWL<3433> A_IWL<3432> A_IWL<3431> A_IWL<3430> A_IWL<3429> A_IWL<3428> A_IWL<3427> A_IWL<3426> A_IWL<3425> A_IWL<3424> A_IWL<3423> A_IWL<3422> A_IWL<3421> A_IWL<3420> A_IWL<3419> A_IWL<3418> A_IWL<3417> A_IWL<3416> A_IWL<3415> A_IWL<3414> A_IWL<3413> A_IWL<3412> A_IWL<3411> A_IWL<3410> A_IWL<3409> A_IWL<3408> A_IWL<3407> A_IWL<3406> A_IWL<3405> A_IWL<3404> A_IWL<3403> A_IWL<3402> A_IWL<3401> A_IWL<3400> A_IWL<3399> A_IWL<3398> A_IWL<3397> A_IWL<3396> A_IWL<3395> A_IWL<3394> A_IWL<3393> A_IWL<3392> A_IWL<3391> A_IWL<3390> A_IWL<3389> A_IWL<3388> A_IWL<3387> A_IWL<3386> A_IWL<3385> A_IWL<3384> A_IWL<3383> A_IWL<3382> A_IWL<3381> A_IWL<3380> A_IWL<3379> A_IWL<3378> A_IWL<3377> A_IWL<3376> A_IWL<3375> A_IWL<3374> A_IWL<3373> A_IWL<3372> A_IWL<3371> A_IWL<3370> A_IWL<3369> A_IWL<3368> A_IWL<3367> A_IWL<3366> A_IWL<3365> A_IWL<3364> A_IWL<3363> A_IWL<3362> A_IWL<3361> A_IWL<3360> A_IWL<3359> A_IWL<3358> A_IWL<3357> A_IWL<3356> A_IWL<3355> A_IWL<3354> A_IWL<3353> A_IWL<3352> A_IWL<3351> A_IWL<3350> A_IWL<3349> A_IWL<3348> A_IWL<3347> A_IWL<3346> A_IWL<3345> A_IWL<3344> A_IWL<3343> A_IWL<3342> A_IWL<3341> A_IWL<3340> A_IWL<3339> A_IWL<3338> A_IWL<3337> A_IWL<3336> A_IWL<3335> A_IWL<3334> A_IWL<3333> A_IWL<3332> A_IWL<3331> A_IWL<3330> A_IWL<3329> A_IWL<3328> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<12> A_BLC<25> A_BLC<24> A_BLC_TOP<25> A_BLC_TOP<24> A_BLT<25> A_BLT<24> A_BLT_TOP<25> A_BLT_TOP<24> A_IWL<3071> A_IWL<3070> A_IWL<3069> A_IWL<3068> A_IWL<3067> A_IWL<3066> A_IWL<3065> A_IWL<3064> A_IWL<3063> A_IWL<3062> A_IWL<3061> A_IWL<3060> A_IWL<3059> A_IWL<3058> A_IWL<3057> A_IWL<3056> A_IWL<3055> A_IWL<3054> A_IWL<3053> A_IWL<3052> A_IWL<3051> A_IWL<3050> A_IWL<3049> A_IWL<3048> A_IWL<3047> A_IWL<3046> A_IWL<3045> A_IWL<3044> A_IWL<3043> A_IWL<3042> A_IWL<3041> A_IWL<3040> A_IWL<3039> A_IWL<3038> A_IWL<3037> A_IWL<3036> A_IWL<3035> A_IWL<3034> A_IWL<3033> A_IWL<3032> A_IWL<3031> A_IWL<3030> A_IWL<3029> A_IWL<3028> A_IWL<3027> A_IWL<3026> A_IWL<3025> A_IWL<3024> A_IWL<3023> A_IWL<3022> A_IWL<3021> A_IWL<3020> A_IWL<3019> A_IWL<3018> A_IWL<3017> A_IWL<3016> A_IWL<3015> A_IWL<3014> A_IWL<3013> A_IWL<3012> A_IWL<3011> A_IWL<3010> A_IWL<3009> A_IWL<3008> A_IWL<3007> A_IWL<3006> A_IWL<3005> A_IWL<3004> A_IWL<3003> A_IWL<3002> A_IWL<3001> A_IWL<3000> A_IWL<2999> A_IWL<2998> A_IWL<2997> A_IWL<2996> A_IWL<2995> A_IWL<2994> A_IWL<2993> A_IWL<2992> A_IWL<2991> A_IWL<2990> A_IWL<2989> A_IWL<2988> A_IWL<2987> A_IWL<2986> A_IWL<2985> A_IWL<2984> A_IWL<2983> A_IWL<2982> A_IWL<2981> A_IWL<2980> A_IWL<2979> A_IWL<2978> A_IWL<2977> A_IWL<2976> A_IWL<2975> A_IWL<2974> A_IWL<2973> A_IWL<2972> A_IWL<2971> A_IWL<2970> A_IWL<2969> A_IWL<2968> A_IWL<2967> A_IWL<2966> A_IWL<2965> A_IWL<2964> A_IWL<2963> A_IWL<2962> A_IWL<2961> A_IWL<2960> A_IWL<2959> A_IWL<2958> A_IWL<2957> A_IWL<2956> A_IWL<2955> A_IWL<2954> A_IWL<2953> A_IWL<2952> A_IWL<2951> A_IWL<2950> A_IWL<2949> A_IWL<2948> A_IWL<2947> A_IWL<2946> A_IWL<2945> A_IWL<2944> A_IWL<2943> A_IWL<2942> A_IWL<2941> A_IWL<2940> A_IWL<2939> A_IWL<2938> A_IWL<2937> A_IWL<2936> A_IWL<2935> A_IWL<2934> A_IWL<2933> A_IWL<2932> A_IWL<2931> A_IWL<2930> A_IWL<2929> A_IWL<2928> A_IWL<2927> A_IWL<2926> A_IWL<2925> A_IWL<2924> A_IWL<2923> A_IWL<2922> A_IWL<2921> A_IWL<2920> A_IWL<2919> A_IWL<2918> A_IWL<2917> A_IWL<2916> A_IWL<2915> A_IWL<2914> A_IWL<2913> A_IWL<2912> A_IWL<2911> A_IWL<2910> A_IWL<2909> A_IWL<2908> A_IWL<2907> A_IWL<2906> A_IWL<2905> A_IWL<2904> A_IWL<2903> A_IWL<2902> A_IWL<2901> A_IWL<2900> A_IWL<2899> A_IWL<2898> A_IWL<2897> A_IWL<2896> A_IWL<2895> A_IWL<2894> A_IWL<2893> A_IWL<2892> A_IWL<2891> A_IWL<2890> A_IWL<2889> A_IWL<2888> A_IWL<2887> A_IWL<2886> A_IWL<2885> A_IWL<2884> A_IWL<2883> A_IWL<2882> A_IWL<2881> A_IWL<2880> A_IWL<2879> A_IWL<2878> A_IWL<2877> A_IWL<2876> A_IWL<2875> A_IWL<2874> A_IWL<2873> A_IWL<2872> A_IWL<2871> A_IWL<2870> A_IWL<2869> A_IWL<2868> A_IWL<2867> A_IWL<2866> A_IWL<2865> A_IWL<2864> A_IWL<2863> A_IWL<2862> A_IWL<2861> A_IWL<2860> A_IWL<2859> A_IWL<2858> A_IWL<2857> A_IWL<2856> A_IWL<2855> A_IWL<2854> A_IWL<2853> A_IWL<2852> A_IWL<2851> A_IWL<2850> A_IWL<2849> A_IWL<2848> A_IWL<2847> A_IWL<2846> A_IWL<2845> A_IWL<2844> A_IWL<2843> A_IWL<2842> A_IWL<2841> A_IWL<2840> A_IWL<2839> A_IWL<2838> A_IWL<2837> A_IWL<2836> A_IWL<2835> A_IWL<2834> A_IWL<2833> A_IWL<2832> A_IWL<2831> A_IWL<2830> A_IWL<2829> A_IWL<2828> A_IWL<2827> A_IWL<2826> A_IWL<2825> A_IWL<2824> A_IWL<2823> A_IWL<2822> A_IWL<2821> A_IWL<2820> A_IWL<2819> A_IWL<2818> A_IWL<2817> A_IWL<2816> A_IWL<3327> A_IWL<3326> A_IWL<3325> A_IWL<3324> A_IWL<3323> A_IWL<3322> A_IWL<3321> A_IWL<3320> A_IWL<3319> A_IWL<3318> A_IWL<3317> A_IWL<3316> A_IWL<3315> A_IWL<3314> A_IWL<3313> A_IWL<3312> A_IWL<3311> A_IWL<3310> A_IWL<3309> A_IWL<3308> A_IWL<3307> A_IWL<3306> A_IWL<3305> A_IWL<3304> A_IWL<3303> A_IWL<3302> A_IWL<3301> A_IWL<3300> A_IWL<3299> A_IWL<3298> A_IWL<3297> A_IWL<3296> A_IWL<3295> A_IWL<3294> A_IWL<3293> A_IWL<3292> A_IWL<3291> A_IWL<3290> A_IWL<3289> A_IWL<3288> A_IWL<3287> A_IWL<3286> A_IWL<3285> A_IWL<3284> A_IWL<3283> A_IWL<3282> A_IWL<3281> A_IWL<3280> A_IWL<3279> A_IWL<3278> A_IWL<3277> A_IWL<3276> A_IWL<3275> A_IWL<3274> A_IWL<3273> A_IWL<3272> A_IWL<3271> A_IWL<3270> A_IWL<3269> A_IWL<3268> A_IWL<3267> A_IWL<3266> A_IWL<3265> A_IWL<3264> A_IWL<3263> A_IWL<3262> A_IWL<3261> A_IWL<3260> A_IWL<3259> A_IWL<3258> A_IWL<3257> A_IWL<3256> A_IWL<3255> A_IWL<3254> A_IWL<3253> A_IWL<3252> A_IWL<3251> A_IWL<3250> A_IWL<3249> A_IWL<3248> A_IWL<3247> A_IWL<3246> A_IWL<3245> A_IWL<3244> A_IWL<3243> A_IWL<3242> A_IWL<3241> A_IWL<3240> A_IWL<3239> A_IWL<3238> A_IWL<3237> A_IWL<3236> A_IWL<3235> A_IWL<3234> A_IWL<3233> A_IWL<3232> A_IWL<3231> A_IWL<3230> A_IWL<3229> A_IWL<3228> A_IWL<3227> A_IWL<3226> A_IWL<3225> A_IWL<3224> A_IWL<3223> A_IWL<3222> A_IWL<3221> A_IWL<3220> A_IWL<3219> A_IWL<3218> A_IWL<3217> A_IWL<3216> A_IWL<3215> A_IWL<3214> A_IWL<3213> A_IWL<3212> A_IWL<3211> A_IWL<3210> A_IWL<3209> A_IWL<3208> A_IWL<3207> A_IWL<3206> A_IWL<3205> A_IWL<3204> A_IWL<3203> A_IWL<3202> A_IWL<3201> A_IWL<3200> A_IWL<3199> A_IWL<3198> A_IWL<3197> A_IWL<3196> A_IWL<3195> A_IWL<3194> A_IWL<3193> A_IWL<3192> A_IWL<3191> A_IWL<3190> A_IWL<3189> A_IWL<3188> A_IWL<3187> A_IWL<3186> A_IWL<3185> A_IWL<3184> A_IWL<3183> A_IWL<3182> A_IWL<3181> A_IWL<3180> A_IWL<3179> A_IWL<3178> A_IWL<3177> A_IWL<3176> A_IWL<3175> A_IWL<3174> A_IWL<3173> A_IWL<3172> A_IWL<3171> A_IWL<3170> A_IWL<3169> A_IWL<3168> A_IWL<3167> A_IWL<3166> A_IWL<3165> A_IWL<3164> A_IWL<3163> A_IWL<3162> A_IWL<3161> A_IWL<3160> A_IWL<3159> A_IWL<3158> A_IWL<3157> A_IWL<3156> A_IWL<3155> A_IWL<3154> A_IWL<3153> A_IWL<3152> A_IWL<3151> A_IWL<3150> A_IWL<3149> A_IWL<3148> A_IWL<3147> A_IWL<3146> A_IWL<3145> A_IWL<3144> A_IWL<3143> A_IWL<3142> A_IWL<3141> A_IWL<3140> A_IWL<3139> A_IWL<3138> A_IWL<3137> A_IWL<3136> A_IWL<3135> A_IWL<3134> A_IWL<3133> A_IWL<3132> A_IWL<3131> A_IWL<3130> A_IWL<3129> A_IWL<3128> A_IWL<3127> A_IWL<3126> A_IWL<3125> A_IWL<3124> A_IWL<3123> A_IWL<3122> A_IWL<3121> A_IWL<3120> A_IWL<3119> A_IWL<3118> A_IWL<3117> A_IWL<3116> A_IWL<3115> A_IWL<3114> A_IWL<3113> A_IWL<3112> A_IWL<3111> A_IWL<3110> A_IWL<3109> A_IWL<3108> A_IWL<3107> A_IWL<3106> A_IWL<3105> A_IWL<3104> A_IWL<3103> A_IWL<3102> A_IWL<3101> A_IWL<3100> A_IWL<3099> A_IWL<3098> A_IWL<3097> A_IWL<3096> A_IWL<3095> A_IWL<3094> A_IWL<3093> A_IWL<3092> A_IWL<3091> A_IWL<3090> A_IWL<3089> A_IWL<3088> A_IWL<3087> A_IWL<3086> A_IWL<3085> A_IWL<3084> A_IWL<3083> A_IWL<3082> A_IWL<3081> A_IWL<3080> A_IWL<3079> A_IWL<3078> A_IWL<3077> A_IWL<3076> A_IWL<3075> A_IWL<3074> A_IWL<3073> A_IWL<3072> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<11> A_BLC<23> A_BLC<22> A_BLC_TOP<23> A_BLC_TOP<22> A_BLT<23> A_BLT<22> A_BLT_TOP<23> A_BLT_TOP<22> A_IWL<2815> A_IWL<2814> A_IWL<2813> A_IWL<2812> A_IWL<2811> A_IWL<2810> A_IWL<2809> A_IWL<2808> A_IWL<2807> A_IWL<2806> A_IWL<2805> A_IWL<2804> A_IWL<2803> A_IWL<2802> A_IWL<2801> A_IWL<2800> A_IWL<2799> A_IWL<2798> A_IWL<2797> A_IWL<2796> A_IWL<2795> A_IWL<2794> A_IWL<2793> A_IWL<2792> A_IWL<2791> A_IWL<2790> A_IWL<2789> A_IWL<2788> A_IWL<2787> A_IWL<2786> A_IWL<2785> A_IWL<2784> A_IWL<2783> A_IWL<2782> A_IWL<2781> A_IWL<2780> A_IWL<2779> A_IWL<2778> A_IWL<2777> A_IWL<2776> A_IWL<2775> A_IWL<2774> A_IWL<2773> A_IWL<2772> A_IWL<2771> A_IWL<2770> A_IWL<2769> A_IWL<2768> A_IWL<2767> A_IWL<2766> A_IWL<2765> A_IWL<2764> A_IWL<2763> A_IWL<2762> A_IWL<2761> A_IWL<2760> A_IWL<2759> A_IWL<2758> A_IWL<2757> A_IWL<2756> A_IWL<2755> A_IWL<2754> A_IWL<2753> A_IWL<2752> A_IWL<2751> A_IWL<2750> A_IWL<2749> A_IWL<2748> A_IWL<2747> A_IWL<2746> A_IWL<2745> A_IWL<2744> A_IWL<2743> A_IWL<2742> A_IWL<2741> A_IWL<2740> A_IWL<2739> A_IWL<2738> A_IWL<2737> A_IWL<2736> A_IWL<2735> A_IWL<2734> A_IWL<2733> A_IWL<2732> A_IWL<2731> A_IWL<2730> A_IWL<2729> A_IWL<2728> A_IWL<2727> A_IWL<2726> A_IWL<2725> A_IWL<2724> A_IWL<2723> A_IWL<2722> A_IWL<2721> A_IWL<2720> A_IWL<2719> A_IWL<2718> A_IWL<2717> A_IWL<2716> A_IWL<2715> A_IWL<2714> A_IWL<2713> A_IWL<2712> A_IWL<2711> A_IWL<2710> A_IWL<2709> A_IWL<2708> A_IWL<2707> A_IWL<2706> A_IWL<2705> A_IWL<2704> A_IWL<2703> A_IWL<2702> A_IWL<2701> A_IWL<2700> A_IWL<2699> A_IWL<2698> A_IWL<2697> A_IWL<2696> A_IWL<2695> A_IWL<2694> A_IWL<2693> A_IWL<2692> A_IWL<2691> A_IWL<2690> A_IWL<2689> A_IWL<2688> A_IWL<2687> A_IWL<2686> A_IWL<2685> A_IWL<2684> A_IWL<2683> A_IWL<2682> A_IWL<2681> A_IWL<2680> A_IWL<2679> A_IWL<2678> A_IWL<2677> A_IWL<2676> A_IWL<2675> A_IWL<2674> A_IWL<2673> A_IWL<2672> A_IWL<2671> A_IWL<2670> A_IWL<2669> A_IWL<2668> A_IWL<2667> A_IWL<2666> A_IWL<2665> A_IWL<2664> A_IWL<2663> A_IWL<2662> A_IWL<2661> A_IWL<2660> A_IWL<2659> A_IWL<2658> A_IWL<2657> A_IWL<2656> A_IWL<2655> A_IWL<2654> A_IWL<2653> A_IWL<2652> A_IWL<2651> A_IWL<2650> A_IWL<2649> A_IWL<2648> A_IWL<2647> A_IWL<2646> A_IWL<2645> A_IWL<2644> A_IWL<2643> A_IWL<2642> A_IWL<2641> A_IWL<2640> A_IWL<2639> A_IWL<2638> A_IWL<2637> A_IWL<2636> A_IWL<2635> A_IWL<2634> A_IWL<2633> A_IWL<2632> A_IWL<2631> A_IWL<2630> A_IWL<2629> A_IWL<2628> A_IWL<2627> A_IWL<2626> A_IWL<2625> A_IWL<2624> A_IWL<2623> A_IWL<2622> A_IWL<2621> A_IWL<2620> A_IWL<2619> A_IWL<2618> A_IWL<2617> A_IWL<2616> A_IWL<2615> A_IWL<2614> A_IWL<2613> A_IWL<2612> A_IWL<2611> A_IWL<2610> A_IWL<2609> A_IWL<2608> A_IWL<2607> A_IWL<2606> A_IWL<2605> A_IWL<2604> A_IWL<2603> A_IWL<2602> A_IWL<2601> A_IWL<2600> A_IWL<2599> A_IWL<2598> A_IWL<2597> A_IWL<2596> A_IWL<2595> A_IWL<2594> A_IWL<2593> A_IWL<2592> A_IWL<2591> A_IWL<2590> A_IWL<2589> A_IWL<2588> A_IWL<2587> A_IWL<2586> A_IWL<2585> A_IWL<2584> A_IWL<2583> A_IWL<2582> A_IWL<2581> A_IWL<2580> A_IWL<2579> A_IWL<2578> A_IWL<2577> A_IWL<2576> A_IWL<2575> A_IWL<2574> A_IWL<2573> A_IWL<2572> A_IWL<2571> A_IWL<2570> A_IWL<2569> A_IWL<2568> A_IWL<2567> A_IWL<2566> A_IWL<2565> A_IWL<2564> A_IWL<2563> A_IWL<2562> A_IWL<2561> A_IWL<2560> A_IWL<3071> A_IWL<3070> A_IWL<3069> A_IWL<3068> A_IWL<3067> A_IWL<3066> A_IWL<3065> A_IWL<3064> A_IWL<3063> A_IWL<3062> A_IWL<3061> A_IWL<3060> A_IWL<3059> A_IWL<3058> A_IWL<3057> A_IWL<3056> A_IWL<3055> A_IWL<3054> A_IWL<3053> A_IWL<3052> A_IWL<3051> A_IWL<3050> A_IWL<3049> A_IWL<3048> A_IWL<3047> A_IWL<3046> A_IWL<3045> A_IWL<3044> A_IWL<3043> A_IWL<3042> A_IWL<3041> A_IWL<3040> A_IWL<3039> A_IWL<3038> A_IWL<3037> A_IWL<3036> A_IWL<3035> A_IWL<3034> A_IWL<3033> A_IWL<3032> A_IWL<3031> A_IWL<3030> A_IWL<3029> A_IWL<3028> A_IWL<3027> A_IWL<3026> A_IWL<3025> A_IWL<3024> A_IWL<3023> A_IWL<3022> A_IWL<3021> A_IWL<3020> A_IWL<3019> A_IWL<3018> A_IWL<3017> A_IWL<3016> A_IWL<3015> A_IWL<3014> A_IWL<3013> A_IWL<3012> A_IWL<3011> A_IWL<3010> A_IWL<3009> A_IWL<3008> A_IWL<3007> A_IWL<3006> A_IWL<3005> A_IWL<3004> A_IWL<3003> A_IWL<3002> A_IWL<3001> A_IWL<3000> A_IWL<2999> A_IWL<2998> A_IWL<2997> A_IWL<2996> A_IWL<2995> A_IWL<2994> A_IWL<2993> A_IWL<2992> A_IWL<2991> A_IWL<2990> A_IWL<2989> A_IWL<2988> A_IWL<2987> A_IWL<2986> A_IWL<2985> A_IWL<2984> A_IWL<2983> A_IWL<2982> A_IWL<2981> A_IWL<2980> A_IWL<2979> A_IWL<2978> A_IWL<2977> A_IWL<2976> A_IWL<2975> A_IWL<2974> A_IWL<2973> A_IWL<2972> A_IWL<2971> A_IWL<2970> A_IWL<2969> A_IWL<2968> A_IWL<2967> A_IWL<2966> A_IWL<2965> A_IWL<2964> A_IWL<2963> A_IWL<2962> A_IWL<2961> A_IWL<2960> A_IWL<2959> A_IWL<2958> A_IWL<2957> A_IWL<2956> A_IWL<2955> A_IWL<2954> A_IWL<2953> A_IWL<2952> A_IWL<2951> A_IWL<2950> A_IWL<2949> A_IWL<2948> A_IWL<2947> A_IWL<2946> A_IWL<2945> A_IWL<2944> A_IWL<2943> A_IWL<2942> A_IWL<2941> A_IWL<2940> A_IWL<2939> A_IWL<2938> A_IWL<2937> A_IWL<2936> A_IWL<2935> A_IWL<2934> A_IWL<2933> A_IWL<2932> A_IWL<2931> A_IWL<2930> A_IWL<2929> A_IWL<2928> A_IWL<2927> A_IWL<2926> A_IWL<2925> A_IWL<2924> A_IWL<2923> A_IWL<2922> A_IWL<2921> A_IWL<2920> A_IWL<2919> A_IWL<2918> A_IWL<2917> A_IWL<2916> A_IWL<2915> A_IWL<2914> A_IWL<2913> A_IWL<2912> A_IWL<2911> A_IWL<2910> A_IWL<2909> A_IWL<2908> A_IWL<2907> A_IWL<2906> A_IWL<2905> A_IWL<2904> A_IWL<2903> A_IWL<2902> A_IWL<2901> A_IWL<2900> A_IWL<2899> A_IWL<2898> A_IWL<2897> A_IWL<2896> A_IWL<2895> A_IWL<2894> A_IWL<2893> A_IWL<2892> A_IWL<2891> A_IWL<2890> A_IWL<2889> A_IWL<2888> A_IWL<2887> A_IWL<2886> A_IWL<2885> A_IWL<2884> A_IWL<2883> A_IWL<2882> A_IWL<2881> A_IWL<2880> A_IWL<2879> A_IWL<2878> A_IWL<2877> A_IWL<2876> A_IWL<2875> A_IWL<2874> A_IWL<2873> A_IWL<2872> A_IWL<2871> A_IWL<2870> A_IWL<2869> A_IWL<2868> A_IWL<2867> A_IWL<2866> A_IWL<2865> A_IWL<2864> A_IWL<2863> A_IWL<2862> A_IWL<2861> A_IWL<2860> A_IWL<2859> A_IWL<2858> A_IWL<2857> A_IWL<2856> A_IWL<2855> A_IWL<2854> A_IWL<2853> A_IWL<2852> A_IWL<2851> A_IWL<2850> A_IWL<2849> A_IWL<2848> A_IWL<2847> A_IWL<2846> A_IWL<2845> A_IWL<2844> A_IWL<2843> A_IWL<2842> A_IWL<2841> A_IWL<2840> A_IWL<2839> A_IWL<2838> A_IWL<2837> A_IWL<2836> A_IWL<2835> A_IWL<2834> A_IWL<2833> A_IWL<2832> A_IWL<2831> A_IWL<2830> A_IWL<2829> A_IWL<2828> A_IWL<2827> A_IWL<2826> A_IWL<2825> A_IWL<2824> A_IWL<2823> A_IWL<2822> A_IWL<2821> A_IWL<2820> A_IWL<2819> A_IWL<2818> A_IWL<2817> A_IWL<2816> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<10> A_BLC<21> A_BLC<20> A_BLC_TOP<21> A_BLC_TOP<20> A_BLT<21> A_BLT<20> A_BLT_TOP<21> A_BLT_TOP<20> A_IWL<2559> A_IWL<2558> A_IWL<2557> A_IWL<2556> A_IWL<2555> A_IWL<2554> A_IWL<2553> A_IWL<2552> A_IWL<2551> A_IWL<2550> A_IWL<2549> A_IWL<2548> A_IWL<2547> A_IWL<2546> A_IWL<2545> A_IWL<2544> A_IWL<2543> A_IWL<2542> A_IWL<2541> A_IWL<2540> A_IWL<2539> A_IWL<2538> A_IWL<2537> A_IWL<2536> A_IWL<2535> A_IWL<2534> A_IWL<2533> A_IWL<2532> A_IWL<2531> A_IWL<2530> A_IWL<2529> A_IWL<2528> A_IWL<2527> A_IWL<2526> A_IWL<2525> A_IWL<2524> A_IWL<2523> A_IWL<2522> A_IWL<2521> A_IWL<2520> A_IWL<2519> A_IWL<2518> A_IWL<2517> A_IWL<2516> A_IWL<2515> A_IWL<2514> A_IWL<2513> A_IWL<2512> A_IWL<2511> A_IWL<2510> A_IWL<2509> A_IWL<2508> A_IWL<2507> A_IWL<2506> A_IWL<2505> A_IWL<2504> A_IWL<2503> A_IWL<2502> A_IWL<2501> A_IWL<2500> A_IWL<2499> A_IWL<2498> A_IWL<2497> A_IWL<2496> A_IWL<2495> A_IWL<2494> A_IWL<2493> A_IWL<2492> A_IWL<2491> A_IWL<2490> A_IWL<2489> A_IWL<2488> A_IWL<2487> A_IWL<2486> A_IWL<2485> A_IWL<2484> A_IWL<2483> A_IWL<2482> A_IWL<2481> A_IWL<2480> A_IWL<2479> A_IWL<2478> A_IWL<2477> A_IWL<2476> A_IWL<2475> A_IWL<2474> A_IWL<2473> A_IWL<2472> A_IWL<2471> A_IWL<2470> A_IWL<2469> A_IWL<2468> A_IWL<2467> A_IWL<2466> A_IWL<2465> A_IWL<2464> A_IWL<2463> A_IWL<2462> A_IWL<2461> A_IWL<2460> A_IWL<2459> A_IWL<2458> A_IWL<2457> A_IWL<2456> A_IWL<2455> A_IWL<2454> A_IWL<2453> A_IWL<2452> A_IWL<2451> A_IWL<2450> A_IWL<2449> A_IWL<2448> A_IWL<2447> A_IWL<2446> A_IWL<2445> A_IWL<2444> A_IWL<2443> A_IWL<2442> A_IWL<2441> A_IWL<2440> A_IWL<2439> A_IWL<2438> A_IWL<2437> A_IWL<2436> A_IWL<2435> A_IWL<2434> A_IWL<2433> A_IWL<2432> A_IWL<2431> A_IWL<2430> A_IWL<2429> A_IWL<2428> A_IWL<2427> A_IWL<2426> A_IWL<2425> A_IWL<2424> A_IWL<2423> A_IWL<2422> A_IWL<2421> A_IWL<2420> A_IWL<2419> A_IWL<2418> A_IWL<2417> A_IWL<2416> A_IWL<2415> A_IWL<2414> A_IWL<2413> A_IWL<2412> A_IWL<2411> A_IWL<2410> A_IWL<2409> A_IWL<2408> A_IWL<2407> A_IWL<2406> A_IWL<2405> A_IWL<2404> A_IWL<2403> A_IWL<2402> A_IWL<2401> A_IWL<2400> A_IWL<2399> A_IWL<2398> A_IWL<2397> A_IWL<2396> A_IWL<2395> A_IWL<2394> A_IWL<2393> A_IWL<2392> A_IWL<2391> A_IWL<2390> A_IWL<2389> A_IWL<2388> A_IWL<2387> A_IWL<2386> A_IWL<2385> A_IWL<2384> A_IWL<2383> A_IWL<2382> A_IWL<2381> A_IWL<2380> A_IWL<2379> A_IWL<2378> A_IWL<2377> A_IWL<2376> A_IWL<2375> A_IWL<2374> A_IWL<2373> A_IWL<2372> A_IWL<2371> A_IWL<2370> A_IWL<2369> A_IWL<2368> A_IWL<2367> A_IWL<2366> A_IWL<2365> A_IWL<2364> A_IWL<2363> A_IWL<2362> A_IWL<2361> A_IWL<2360> A_IWL<2359> A_IWL<2358> A_IWL<2357> A_IWL<2356> A_IWL<2355> A_IWL<2354> A_IWL<2353> A_IWL<2352> A_IWL<2351> A_IWL<2350> A_IWL<2349> A_IWL<2348> A_IWL<2347> A_IWL<2346> A_IWL<2345> A_IWL<2344> A_IWL<2343> A_IWL<2342> A_IWL<2341> A_IWL<2340> A_IWL<2339> A_IWL<2338> A_IWL<2337> A_IWL<2336> A_IWL<2335> A_IWL<2334> A_IWL<2333> A_IWL<2332> A_IWL<2331> A_IWL<2330> A_IWL<2329> A_IWL<2328> A_IWL<2327> A_IWL<2326> A_IWL<2325> A_IWL<2324> A_IWL<2323> A_IWL<2322> A_IWL<2321> A_IWL<2320> A_IWL<2319> A_IWL<2318> A_IWL<2317> A_IWL<2316> A_IWL<2315> A_IWL<2314> A_IWL<2313> A_IWL<2312> A_IWL<2311> A_IWL<2310> A_IWL<2309> A_IWL<2308> A_IWL<2307> A_IWL<2306> A_IWL<2305> A_IWL<2304> A_IWL<2815> A_IWL<2814> A_IWL<2813> A_IWL<2812> A_IWL<2811> A_IWL<2810> A_IWL<2809> A_IWL<2808> A_IWL<2807> A_IWL<2806> A_IWL<2805> A_IWL<2804> A_IWL<2803> A_IWL<2802> A_IWL<2801> A_IWL<2800> A_IWL<2799> A_IWL<2798> A_IWL<2797> A_IWL<2796> A_IWL<2795> A_IWL<2794> A_IWL<2793> A_IWL<2792> A_IWL<2791> A_IWL<2790> A_IWL<2789> A_IWL<2788> A_IWL<2787> A_IWL<2786> A_IWL<2785> A_IWL<2784> A_IWL<2783> A_IWL<2782> A_IWL<2781> A_IWL<2780> A_IWL<2779> A_IWL<2778> A_IWL<2777> A_IWL<2776> A_IWL<2775> A_IWL<2774> A_IWL<2773> A_IWL<2772> A_IWL<2771> A_IWL<2770> A_IWL<2769> A_IWL<2768> A_IWL<2767> A_IWL<2766> A_IWL<2765> A_IWL<2764> A_IWL<2763> A_IWL<2762> A_IWL<2761> A_IWL<2760> A_IWL<2759> A_IWL<2758> A_IWL<2757> A_IWL<2756> A_IWL<2755> A_IWL<2754> A_IWL<2753> A_IWL<2752> A_IWL<2751> A_IWL<2750> A_IWL<2749> A_IWL<2748> A_IWL<2747> A_IWL<2746> A_IWL<2745> A_IWL<2744> A_IWL<2743> A_IWL<2742> A_IWL<2741> A_IWL<2740> A_IWL<2739> A_IWL<2738> A_IWL<2737> A_IWL<2736> A_IWL<2735> A_IWL<2734> A_IWL<2733> A_IWL<2732> A_IWL<2731> A_IWL<2730> A_IWL<2729> A_IWL<2728> A_IWL<2727> A_IWL<2726> A_IWL<2725> A_IWL<2724> A_IWL<2723> A_IWL<2722> A_IWL<2721> A_IWL<2720> A_IWL<2719> A_IWL<2718> A_IWL<2717> A_IWL<2716> A_IWL<2715> A_IWL<2714> A_IWL<2713> A_IWL<2712> A_IWL<2711> A_IWL<2710> A_IWL<2709> A_IWL<2708> A_IWL<2707> A_IWL<2706> A_IWL<2705> A_IWL<2704> A_IWL<2703> A_IWL<2702> A_IWL<2701> A_IWL<2700> A_IWL<2699> A_IWL<2698> A_IWL<2697> A_IWL<2696> A_IWL<2695> A_IWL<2694> A_IWL<2693> A_IWL<2692> A_IWL<2691> A_IWL<2690> A_IWL<2689> A_IWL<2688> A_IWL<2687> A_IWL<2686> A_IWL<2685> A_IWL<2684> A_IWL<2683> A_IWL<2682> A_IWL<2681> A_IWL<2680> A_IWL<2679> A_IWL<2678> A_IWL<2677> A_IWL<2676> A_IWL<2675> A_IWL<2674> A_IWL<2673> A_IWL<2672> A_IWL<2671> A_IWL<2670> A_IWL<2669> A_IWL<2668> A_IWL<2667> A_IWL<2666> A_IWL<2665> A_IWL<2664> A_IWL<2663> A_IWL<2662> A_IWL<2661> A_IWL<2660> A_IWL<2659> A_IWL<2658> A_IWL<2657> A_IWL<2656> A_IWL<2655> A_IWL<2654> A_IWL<2653> A_IWL<2652> A_IWL<2651> A_IWL<2650> A_IWL<2649> A_IWL<2648> A_IWL<2647> A_IWL<2646> A_IWL<2645> A_IWL<2644> A_IWL<2643> A_IWL<2642> A_IWL<2641> A_IWL<2640> A_IWL<2639> A_IWL<2638> A_IWL<2637> A_IWL<2636> A_IWL<2635> A_IWL<2634> A_IWL<2633> A_IWL<2632> A_IWL<2631> A_IWL<2630> A_IWL<2629> A_IWL<2628> A_IWL<2627> A_IWL<2626> A_IWL<2625> A_IWL<2624> A_IWL<2623> A_IWL<2622> A_IWL<2621> A_IWL<2620> A_IWL<2619> A_IWL<2618> A_IWL<2617> A_IWL<2616> A_IWL<2615> A_IWL<2614> A_IWL<2613> A_IWL<2612> A_IWL<2611> A_IWL<2610> A_IWL<2609> A_IWL<2608> A_IWL<2607> A_IWL<2606> A_IWL<2605> A_IWL<2604> A_IWL<2603> A_IWL<2602> A_IWL<2601> A_IWL<2600> A_IWL<2599> A_IWL<2598> A_IWL<2597> A_IWL<2596> A_IWL<2595> A_IWL<2594> A_IWL<2593> A_IWL<2592> A_IWL<2591> A_IWL<2590> A_IWL<2589> A_IWL<2588> A_IWL<2587> A_IWL<2586> A_IWL<2585> A_IWL<2584> A_IWL<2583> A_IWL<2582> A_IWL<2581> A_IWL<2580> A_IWL<2579> A_IWL<2578> A_IWL<2577> A_IWL<2576> A_IWL<2575> A_IWL<2574> A_IWL<2573> A_IWL<2572> A_IWL<2571> A_IWL<2570> A_IWL<2569> A_IWL<2568> A_IWL<2567> A_IWL<2566> A_IWL<2565> A_IWL<2564> A_IWL<2563> A_IWL<2562> A_IWL<2561> A_IWL<2560> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<9> A_BLC<19> A_BLC<18> A_BLC_TOP<19> A_BLC_TOP<18> A_BLT<19> A_BLT<18> A_BLT_TOP<19> A_BLT_TOP<18> A_IWL<2303> A_IWL<2302> A_IWL<2301> A_IWL<2300> A_IWL<2299> A_IWL<2298> A_IWL<2297> A_IWL<2296> A_IWL<2295> A_IWL<2294> A_IWL<2293> A_IWL<2292> A_IWL<2291> A_IWL<2290> A_IWL<2289> A_IWL<2288> A_IWL<2287> A_IWL<2286> A_IWL<2285> A_IWL<2284> A_IWL<2283> A_IWL<2282> A_IWL<2281> A_IWL<2280> A_IWL<2279> A_IWL<2278> A_IWL<2277> A_IWL<2276> A_IWL<2275> A_IWL<2274> A_IWL<2273> A_IWL<2272> A_IWL<2271> A_IWL<2270> A_IWL<2269> A_IWL<2268> A_IWL<2267> A_IWL<2266> A_IWL<2265> A_IWL<2264> A_IWL<2263> A_IWL<2262> A_IWL<2261> A_IWL<2260> A_IWL<2259> A_IWL<2258> A_IWL<2257> A_IWL<2256> A_IWL<2255> A_IWL<2254> A_IWL<2253> A_IWL<2252> A_IWL<2251> A_IWL<2250> A_IWL<2249> A_IWL<2248> A_IWL<2247> A_IWL<2246> A_IWL<2245> A_IWL<2244> A_IWL<2243> A_IWL<2242> A_IWL<2241> A_IWL<2240> A_IWL<2239> A_IWL<2238> A_IWL<2237> A_IWL<2236> A_IWL<2235> A_IWL<2234> A_IWL<2233> A_IWL<2232> A_IWL<2231> A_IWL<2230> A_IWL<2229> A_IWL<2228> A_IWL<2227> A_IWL<2226> A_IWL<2225> A_IWL<2224> A_IWL<2223> A_IWL<2222> A_IWL<2221> A_IWL<2220> A_IWL<2219> A_IWL<2218> A_IWL<2217> A_IWL<2216> A_IWL<2215> A_IWL<2214> A_IWL<2213> A_IWL<2212> A_IWL<2211> A_IWL<2210> A_IWL<2209> A_IWL<2208> A_IWL<2207> A_IWL<2206> A_IWL<2205> A_IWL<2204> A_IWL<2203> A_IWL<2202> A_IWL<2201> A_IWL<2200> A_IWL<2199> A_IWL<2198> A_IWL<2197> A_IWL<2196> A_IWL<2195> A_IWL<2194> A_IWL<2193> A_IWL<2192> A_IWL<2191> A_IWL<2190> A_IWL<2189> A_IWL<2188> A_IWL<2187> A_IWL<2186> A_IWL<2185> A_IWL<2184> A_IWL<2183> A_IWL<2182> A_IWL<2181> A_IWL<2180> A_IWL<2179> A_IWL<2178> A_IWL<2177> A_IWL<2176> A_IWL<2175> A_IWL<2174> A_IWL<2173> A_IWL<2172> A_IWL<2171> A_IWL<2170> A_IWL<2169> A_IWL<2168> A_IWL<2167> A_IWL<2166> A_IWL<2165> A_IWL<2164> A_IWL<2163> A_IWL<2162> A_IWL<2161> A_IWL<2160> A_IWL<2159> A_IWL<2158> A_IWL<2157> A_IWL<2156> A_IWL<2155> A_IWL<2154> A_IWL<2153> A_IWL<2152> A_IWL<2151> A_IWL<2150> A_IWL<2149> A_IWL<2148> A_IWL<2147> A_IWL<2146> A_IWL<2145> A_IWL<2144> A_IWL<2143> A_IWL<2142> A_IWL<2141> A_IWL<2140> A_IWL<2139> A_IWL<2138> A_IWL<2137> A_IWL<2136> A_IWL<2135> A_IWL<2134> A_IWL<2133> A_IWL<2132> A_IWL<2131> A_IWL<2130> A_IWL<2129> A_IWL<2128> A_IWL<2127> A_IWL<2126> A_IWL<2125> A_IWL<2124> A_IWL<2123> A_IWL<2122> A_IWL<2121> A_IWL<2120> A_IWL<2119> A_IWL<2118> A_IWL<2117> A_IWL<2116> A_IWL<2115> A_IWL<2114> A_IWL<2113> A_IWL<2112> A_IWL<2111> A_IWL<2110> A_IWL<2109> A_IWL<2108> A_IWL<2107> A_IWL<2106> A_IWL<2105> A_IWL<2104> A_IWL<2103> A_IWL<2102> A_IWL<2101> A_IWL<2100> A_IWL<2099> A_IWL<2098> A_IWL<2097> A_IWL<2096> A_IWL<2095> A_IWL<2094> A_IWL<2093> A_IWL<2092> A_IWL<2091> A_IWL<2090> A_IWL<2089> A_IWL<2088> A_IWL<2087> A_IWL<2086> A_IWL<2085> A_IWL<2084> A_IWL<2083> A_IWL<2082> A_IWL<2081> A_IWL<2080> A_IWL<2079> A_IWL<2078> A_IWL<2077> A_IWL<2076> A_IWL<2075> A_IWL<2074> A_IWL<2073> A_IWL<2072> A_IWL<2071> A_IWL<2070> A_IWL<2069> A_IWL<2068> A_IWL<2067> A_IWL<2066> A_IWL<2065> A_IWL<2064> A_IWL<2063> A_IWL<2062> A_IWL<2061> A_IWL<2060> A_IWL<2059> A_IWL<2058> A_IWL<2057> A_IWL<2056> A_IWL<2055> A_IWL<2054> A_IWL<2053> A_IWL<2052> A_IWL<2051> A_IWL<2050> A_IWL<2049> A_IWL<2048> A_IWL<2559> A_IWL<2558> A_IWL<2557> A_IWL<2556> A_IWL<2555> A_IWL<2554> A_IWL<2553> A_IWL<2552> A_IWL<2551> A_IWL<2550> A_IWL<2549> A_IWL<2548> A_IWL<2547> A_IWL<2546> A_IWL<2545> A_IWL<2544> A_IWL<2543> A_IWL<2542> A_IWL<2541> A_IWL<2540> A_IWL<2539> A_IWL<2538> A_IWL<2537> A_IWL<2536> A_IWL<2535> A_IWL<2534> A_IWL<2533> A_IWL<2532> A_IWL<2531> A_IWL<2530> A_IWL<2529> A_IWL<2528> A_IWL<2527> A_IWL<2526> A_IWL<2525> A_IWL<2524> A_IWL<2523> A_IWL<2522> A_IWL<2521> A_IWL<2520> A_IWL<2519> A_IWL<2518> A_IWL<2517> A_IWL<2516> A_IWL<2515> A_IWL<2514> A_IWL<2513> A_IWL<2512> A_IWL<2511> A_IWL<2510> A_IWL<2509> A_IWL<2508> A_IWL<2507> A_IWL<2506> A_IWL<2505> A_IWL<2504> A_IWL<2503> A_IWL<2502> A_IWL<2501> A_IWL<2500> A_IWL<2499> A_IWL<2498> A_IWL<2497> A_IWL<2496> A_IWL<2495> A_IWL<2494> A_IWL<2493> A_IWL<2492> A_IWL<2491> A_IWL<2490> A_IWL<2489> A_IWL<2488> A_IWL<2487> A_IWL<2486> A_IWL<2485> A_IWL<2484> A_IWL<2483> A_IWL<2482> A_IWL<2481> A_IWL<2480> A_IWL<2479> A_IWL<2478> A_IWL<2477> A_IWL<2476> A_IWL<2475> A_IWL<2474> A_IWL<2473> A_IWL<2472> A_IWL<2471> A_IWL<2470> A_IWL<2469> A_IWL<2468> A_IWL<2467> A_IWL<2466> A_IWL<2465> A_IWL<2464> A_IWL<2463> A_IWL<2462> A_IWL<2461> A_IWL<2460> A_IWL<2459> A_IWL<2458> A_IWL<2457> A_IWL<2456> A_IWL<2455> A_IWL<2454> A_IWL<2453> A_IWL<2452> A_IWL<2451> A_IWL<2450> A_IWL<2449> A_IWL<2448> A_IWL<2447> A_IWL<2446> A_IWL<2445> A_IWL<2444> A_IWL<2443> A_IWL<2442> A_IWL<2441> A_IWL<2440> A_IWL<2439> A_IWL<2438> A_IWL<2437> A_IWL<2436> A_IWL<2435> A_IWL<2434> A_IWL<2433> A_IWL<2432> A_IWL<2431> A_IWL<2430> A_IWL<2429> A_IWL<2428> A_IWL<2427> A_IWL<2426> A_IWL<2425> A_IWL<2424> A_IWL<2423> A_IWL<2422> A_IWL<2421> A_IWL<2420> A_IWL<2419> A_IWL<2418> A_IWL<2417> A_IWL<2416> A_IWL<2415> A_IWL<2414> A_IWL<2413> A_IWL<2412> A_IWL<2411> A_IWL<2410> A_IWL<2409> A_IWL<2408> A_IWL<2407> A_IWL<2406> A_IWL<2405> A_IWL<2404> A_IWL<2403> A_IWL<2402> A_IWL<2401> A_IWL<2400> A_IWL<2399> A_IWL<2398> A_IWL<2397> A_IWL<2396> A_IWL<2395> A_IWL<2394> A_IWL<2393> A_IWL<2392> A_IWL<2391> A_IWL<2390> A_IWL<2389> A_IWL<2388> A_IWL<2387> A_IWL<2386> A_IWL<2385> A_IWL<2384> A_IWL<2383> A_IWL<2382> A_IWL<2381> A_IWL<2380> A_IWL<2379> A_IWL<2378> A_IWL<2377> A_IWL<2376> A_IWL<2375> A_IWL<2374> A_IWL<2373> A_IWL<2372> A_IWL<2371> A_IWL<2370> A_IWL<2369> A_IWL<2368> A_IWL<2367> A_IWL<2366> A_IWL<2365> A_IWL<2364> A_IWL<2363> A_IWL<2362> A_IWL<2361> A_IWL<2360> A_IWL<2359> A_IWL<2358> A_IWL<2357> A_IWL<2356> A_IWL<2355> A_IWL<2354> A_IWL<2353> A_IWL<2352> A_IWL<2351> A_IWL<2350> A_IWL<2349> A_IWL<2348> A_IWL<2347> A_IWL<2346> A_IWL<2345> A_IWL<2344> A_IWL<2343> A_IWL<2342> A_IWL<2341> A_IWL<2340> A_IWL<2339> A_IWL<2338> A_IWL<2337> A_IWL<2336> A_IWL<2335> A_IWL<2334> A_IWL<2333> A_IWL<2332> A_IWL<2331> A_IWL<2330> A_IWL<2329> A_IWL<2328> A_IWL<2327> A_IWL<2326> A_IWL<2325> A_IWL<2324> A_IWL<2323> A_IWL<2322> A_IWL<2321> A_IWL<2320> A_IWL<2319> A_IWL<2318> A_IWL<2317> A_IWL<2316> A_IWL<2315> A_IWL<2314> A_IWL<2313> A_IWL<2312> A_IWL<2311> A_IWL<2310> A_IWL<2309> A_IWL<2308> A_IWL<2307> A_IWL<2306> A_IWL<2305> A_IWL<2304> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<8> A_BLC<17> A_BLC<16> A_BLC_TOP<17> A_BLC_TOP<16> A_BLT<17> A_BLT<16> A_BLT_TOP<17> A_BLT_TOP<16> A_IWL<2047> A_IWL<2046> A_IWL<2045> A_IWL<2044> A_IWL<2043> A_IWL<2042> A_IWL<2041> A_IWL<2040> A_IWL<2039> A_IWL<2038> A_IWL<2037> A_IWL<2036> A_IWL<2035> A_IWL<2034> A_IWL<2033> A_IWL<2032> A_IWL<2031> A_IWL<2030> A_IWL<2029> A_IWL<2028> A_IWL<2027> A_IWL<2026> A_IWL<2025> A_IWL<2024> A_IWL<2023> A_IWL<2022> A_IWL<2021> A_IWL<2020> A_IWL<2019> A_IWL<2018> A_IWL<2017> A_IWL<2016> A_IWL<2015> A_IWL<2014> A_IWL<2013> A_IWL<2012> A_IWL<2011> A_IWL<2010> A_IWL<2009> A_IWL<2008> A_IWL<2007> A_IWL<2006> A_IWL<2005> A_IWL<2004> A_IWL<2003> A_IWL<2002> A_IWL<2001> A_IWL<2000> A_IWL<1999> A_IWL<1998> A_IWL<1997> A_IWL<1996> A_IWL<1995> A_IWL<1994> A_IWL<1993> A_IWL<1992> A_IWL<1991> A_IWL<1990> A_IWL<1989> A_IWL<1988> A_IWL<1987> A_IWL<1986> A_IWL<1985> A_IWL<1984> A_IWL<1983> A_IWL<1982> A_IWL<1981> A_IWL<1980> A_IWL<1979> A_IWL<1978> A_IWL<1977> A_IWL<1976> A_IWL<1975> A_IWL<1974> A_IWL<1973> A_IWL<1972> A_IWL<1971> A_IWL<1970> A_IWL<1969> A_IWL<1968> A_IWL<1967> A_IWL<1966> A_IWL<1965> A_IWL<1964> A_IWL<1963> A_IWL<1962> A_IWL<1961> A_IWL<1960> A_IWL<1959> A_IWL<1958> A_IWL<1957> A_IWL<1956> A_IWL<1955> A_IWL<1954> A_IWL<1953> A_IWL<1952> A_IWL<1951> A_IWL<1950> A_IWL<1949> A_IWL<1948> A_IWL<1947> A_IWL<1946> A_IWL<1945> A_IWL<1944> A_IWL<1943> A_IWL<1942> A_IWL<1941> A_IWL<1940> A_IWL<1939> A_IWL<1938> A_IWL<1937> A_IWL<1936> A_IWL<1935> A_IWL<1934> A_IWL<1933> A_IWL<1932> A_IWL<1931> A_IWL<1930> A_IWL<1929> A_IWL<1928> A_IWL<1927> A_IWL<1926> A_IWL<1925> A_IWL<1924> A_IWL<1923> A_IWL<1922> A_IWL<1921> A_IWL<1920> A_IWL<1919> A_IWL<1918> A_IWL<1917> A_IWL<1916> A_IWL<1915> A_IWL<1914> A_IWL<1913> A_IWL<1912> A_IWL<1911> A_IWL<1910> A_IWL<1909> A_IWL<1908> A_IWL<1907> A_IWL<1906> A_IWL<1905> A_IWL<1904> A_IWL<1903> A_IWL<1902> A_IWL<1901> A_IWL<1900> A_IWL<1899> A_IWL<1898> A_IWL<1897> A_IWL<1896> A_IWL<1895> A_IWL<1894> A_IWL<1893> A_IWL<1892> A_IWL<1891> A_IWL<1890> A_IWL<1889> A_IWL<1888> A_IWL<1887> A_IWL<1886> A_IWL<1885> A_IWL<1884> A_IWL<1883> A_IWL<1882> A_IWL<1881> A_IWL<1880> A_IWL<1879> A_IWL<1878> A_IWL<1877> A_IWL<1876> A_IWL<1875> A_IWL<1874> A_IWL<1873> A_IWL<1872> A_IWL<1871> A_IWL<1870> A_IWL<1869> A_IWL<1868> A_IWL<1867> A_IWL<1866> A_IWL<1865> A_IWL<1864> A_IWL<1863> A_IWL<1862> A_IWL<1861> A_IWL<1860> A_IWL<1859> A_IWL<1858> A_IWL<1857> A_IWL<1856> A_IWL<1855> A_IWL<1854> A_IWL<1853> A_IWL<1852> A_IWL<1851> A_IWL<1850> A_IWL<1849> A_IWL<1848> A_IWL<1847> A_IWL<1846> A_IWL<1845> A_IWL<1844> A_IWL<1843> A_IWL<1842> A_IWL<1841> A_IWL<1840> A_IWL<1839> A_IWL<1838> A_IWL<1837> A_IWL<1836> A_IWL<1835> A_IWL<1834> A_IWL<1833> A_IWL<1832> A_IWL<1831> A_IWL<1830> A_IWL<1829> A_IWL<1828> A_IWL<1827> A_IWL<1826> A_IWL<1825> A_IWL<1824> A_IWL<1823> A_IWL<1822> A_IWL<1821> A_IWL<1820> A_IWL<1819> A_IWL<1818> A_IWL<1817> A_IWL<1816> A_IWL<1815> A_IWL<1814> A_IWL<1813> A_IWL<1812> A_IWL<1811> A_IWL<1810> A_IWL<1809> A_IWL<1808> A_IWL<1807> A_IWL<1806> A_IWL<1805> A_IWL<1804> A_IWL<1803> A_IWL<1802> A_IWL<1801> A_IWL<1800> A_IWL<1799> A_IWL<1798> A_IWL<1797> A_IWL<1796> A_IWL<1795> A_IWL<1794> A_IWL<1793> A_IWL<1792> A_IWL<2303> A_IWL<2302> A_IWL<2301> A_IWL<2300> A_IWL<2299> A_IWL<2298> A_IWL<2297> A_IWL<2296> A_IWL<2295> A_IWL<2294> A_IWL<2293> A_IWL<2292> A_IWL<2291> A_IWL<2290> A_IWL<2289> A_IWL<2288> A_IWL<2287> A_IWL<2286> A_IWL<2285> A_IWL<2284> A_IWL<2283> A_IWL<2282> A_IWL<2281> A_IWL<2280> A_IWL<2279> A_IWL<2278> A_IWL<2277> A_IWL<2276> A_IWL<2275> A_IWL<2274> A_IWL<2273> A_IWL<2272> A_IWL<2271> A_IWL<2270> A_IWL<2269> A_IWL<2268> A_IWL<2267> A_IWL<2266> A_IWL<2265> A_IWL<2264> A_IWL<2263> A_IWL<2262> A_IWL<2261> A_IWL<2260> A_IWL<2259> A_IWL<2258> A_IWL<2257> A_IWL<2256> A_IWL<2255> A_IWL<2254> A_IWL<2253> A_IWL<2252> A_IWL<2251> A_IWL<2250> A_IWL<2249> A_IWL<2248> A_IWL<2247> A_IWL<2246> A_IWL<2245> A_IWL<2244> A_IWL<2243> A_IWL<2242> A_IWL<2241> A_IWL<2240> A_IWL<2239> A_IWL<2238> A_IWL<2237> A_IWL<2236> A_IWL<2235> A_IWL<2234> A_IWL<2233> A_IWL<2232> A_IWL<2231> A_IWL<2230> A_IWL<2229> A_IWL<2228> A_IWL<2227> A_IWL<2226> A_IWL<2225> A_IWL<2224> A_IWL<2223> A_IWL<2222> A_IWL<2221> A_IWL<2220> A_IWL<2219> A_IWL<2218> A_IWL<2217> A_IWL<2216> A_IWL<2215> A_IWL<2214> A_IWL<2213> A_IWL<2212> A_IWL<2211> A_IWL<2210> A_IWL<2209> A_IWL<2208> A_IWL<2207> A_IWL<2206> A_IWL<2205> A_IWL<2204> A_IWL<2203> A_IWL<2202> A_IWL<2201> A_IWL<2200> A_IWL<2199> A_IWL<2198> A_IWL<2197> A_IWL<2196> A_IWL<2195> A_IWL<2194> A_IWL<2193> A_IWL<2192> A_IWL<2191> A_IWL<2190> A_IWL<2189> A_IWL<2188> A_IWL<2187> A_IWL<2186> A_IWL<2185> A_IWL<2184> A_IWL<2183> A_IWL<2182> A_IWL<2181> A_IWL<2180> A_IWL<2179> A_IWL<2178> A_IWL<2177> A_IWL<2176> A_IWL<2175> A_IWL<2174> A_IWL<2173> A_IWL<2172> A_IWL<2171> A_IWL<2170> A_IWL<2169> A_IWL<2168> A_IWL<2167> A_IWL<2166> A_IWL<2165> A_IWL<2164> A_IWL<2163> A_IWL<2162> A_IWL<2161> A_IWL<2160> A_IWL<2159> A_IWL<2158> A_IWL<2157> A_IWL<2156> A_IWL<2155> A_IWL<2154> A_IWL<2153> A_IWL<2152> A_IWL<2151> A_IWL<2150> A_IWL<2149> A_IWL<2148> A_IWL<2147> A_IWL<2146> A_IWL<2145> A_IWL<2144> A_IWL<2143> A_IWL<2142> A_IWL<2141> A_IWL<2140> A_IWL<2139> A_IWL<2138> A_IWL<2137> A_IWL<2136> A_IWL<2135> A_IWL<2134> A_IWL<2133> A_IWL<2132> A_IWL<2131> A_IWL<2130> A_IWL<2129> A_IWL<2128> A_IWL<2127> A_IWL<2126> A_IWL<2125> A_IWL<2124> A_IWL<2123> A_IWL<2122> A_IWL<2121> A_IWL<2120> A_IWL<2119> A_IWL<2118> A_IWL<2117> A_IWL<2116> A_IWL<2115> A_IWL<2114> A_IWL<2113> A_IWL<2112> A_IWL<2111> A_IWL<2110> A_IWL<2109> A_IWL<2108> A_IWL<2107> A_IWL<2106> A_IWL<2105> A_IWL<2104> A_IWL<2103> A_IWL<2102> A_IWL<2101> A_IWL<2100> A_IWL<2099> A_IWL<2098> A_IWL<2097> A_IWL<2096> A_IWL<2095> A_IWL<2094> A_IWL<2093> A_IWL<2092> A_IWL<2091> A_IWL<2090> A_IWL<2089> A_IWL<2088> A_IWL<2087> A_IWL<2086> A_IWL<2085> A_IWL<2084> A_IWL<2083> A_IWL<2082> A_IWL<2081> A_IWL<2080> A_IWL<2079> A_IWL<2078> A_IWL<2077> A_IWL<2076> A_IWL<2075> A_IWL<2074> A_IWL<2073> A_IWL<2072> A_IWL<2071> A_IWL<2070> A_IWL<2069> A_IWL<2068> A_IWL<2067> A_IWL<2066> A_IWL<2065> A_IWL<2064> A_IWL<2063> A_IWL<2062> A_IWL<2061> A_IWL<2060> A_IWL<2059> A_IWL<2058> A_IWL<2057> A_IWL<2056> A_IWL<2055> A_IWL<2054> A_IWL<2053> A_IWL<2052> A_IWL<2051> A_IWL<2050> A_IWL<2049> A_IWL<2048> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<7> A_BLC<15> A_BLC<14> A_BLC_TOP<15> A_BLC_TOP<14> A_BLT<15> A_BLT<14> A_BLT_TOP<15> A_BLT_TOP<14> A_IWL<1791> A_IWL<1790> A_IWL<1789> A_IWL<1788> A_IWL<1787> A_IWL<1786> A_IWL<1785> A_IWL<1784> A_IWL<1783> A_IWL<1782> A_IWL<1781> A_IWL<1780> A_IWL<1779> A_IWL<1778> A_IWL<1777> A_IWL<1776> A_IWL<1775> A_IWL<1774> A_IWL<1773> A_IWL<1772> A_IWL<1771> A_IWL<1770> A_IWL<1769> A_IWL<1768> A_IWL<1767> A_IWL<1766> A_IWL<1765> A_IWL<1764> A_IWL<1763> A_IWL<1762> A_IWL<1761> A_IWL<1760> A_IWL<1759> A_IWL<1758> A_IWL<1757> A_IWL<1756> A_IWL<1755> A_IWL<1754> A_IWL<1753> A_IWL<1752> A_IWL<1751> A_IWL<1750> A_IWL<1749> A_IWL<1748> A_IWL<1747> A_IWL<1746> A_IWL<1745> A_IWL<1744> A_IWL<1743> A_IWL<1742> A_IWL<1741> A_IWL<1740> A_IWL<1739> A_IWL<1738> A_IWL<1737> A_IWL<1736> A_IWL<1735> A_IWL<1734> A_IWL<1733> A_IWL<1732> A_IWL<1731> A_IWL<1730> A_IWL<1729> A_IWL<1728> A_IWL<1727> A_IWL<1726> A_IWL<1725> A_IWL<1724> A_IWL<1723> A_IWL<1722> A_IWL<1721> A_IWL<1720> A_IWL<1719> A_IWL<1718> A_IWL<1717> A_IWL<1716> A_IWL<1715> A_IWL<1714> A_IWL<1713> A_IWL<1712> A_IWL<1711> A_IWL<1710> A_IWL<1709> A_IWL<1708> A_IWL<1707> A_IWL<1706> A_IWL<1705> A_IWL<1704> A_IWL<1703> A_IWL<1702> A_IWL<1701> A_IWL<1700> A_IWL<1699> A_IWL<1698> A_IWL<1697> A_IWL<1696> A_IWL<1695> A_IWL<1694> A_IWL<1693> A_IWL<1692> A_IWL<1691> A_IWL<1690> A_IWL<1689> A_IWL<1688> A_IWL<1687> A_IWL<1686> A_IWL<1685> A_IWL<1684> A_IWL<1683> A_IWL<1682> A_IWL<1681> A_IWL<1680> A_IWL<1679> A_IWL<1678> A_IWL<1677> A_IWL<1676> A_IWL<1675> A_IWL<1674> A_IWL<1673> A_IWL<1672> A_IWL<1671> A_IWL<1670> A_IWL<1669> A_IWL<1668> A_IWL<1667> A_IWL<1666> A_IWL<1665> A_IWL<1664> A_IWL<1663> A_IWL<1662> A_IWL<1661> A_IWL<1660> A_IWL<1659> A_IWL<1658> A_IWL<1657> A_IWL<1656> A_IWL<1655> A_IWL<1654> A_IWL<1653> A_IWL<1652> A_IWL<1651> A_IWL<1650> A_IWL<1649> A_IWL<1648> A_IWL<1647> A_IWL<1646> A_IWL<1645> A_IWL<1644> A_IWL<1643> A_IWL<1642> A_IWL<1641> A_IWL<1640> A_IWL<1639> A_IWL<1638> A_IWL<1637> A_IWL<1636> A_IWL<1635> A_IWL<1634> A_IWL<1633> A_IWL<1632> A_IWL<1631> A_IWL<1630> A_IWL<1629> A_IWL<1628> A_IWL<1627> A_IWL<1626> A_IWL<1625> A_IWL<1624> A_IWL<1623> A_IWL<1622> A_IWL<1621> A_IWL<1620> A_IWL<1619> A_IWL<1618> A_IWL<1617> A_IWL<1616> A_IWL<1615> A_IWL<1614> A_IWL<1613> A_IWL<1612> A_IWL<1611> A_IWL<1610> A_IWL<1609> A_IWL<1608> A_IWL<1607> A_IWL<1606> A_IWL<1605> A_IWL<1604> A_IWL<1603> A_IWL<1602> A_IWL<1601> A_IWL<1600> A_IWL<1599> A_IWL<1598> A_IWL<1597> A_IWL<1596> A_IWL<1595> A_IWL<1594> A_IWL<1593> A_IWL<1592> A_IWL<1591> A_IWL<1590> A_IWL<1589> A_IWL<1588> A_IWL<1587> A_IWL<1586> A_IWL<1585> A_IWL<1584> A_IWL<1583> A_IWL<1582> A_IWL<1581> A_IWL<1580> A_IWL<1579> A_IWL<1578> A_IWL<1577> A_IWL<1576> A_IWL<1575> A_IWL<1574> A_IWL<1573> A_IWL<1572> A_IWL<1571> A_IWL<1570> A_IWL<1569> A_IWL<1568> A_IWL<1567> A_IWL<1566> A_IWL<1565> A_IWL<1564> A_IWL<1563> A_IWL<1562> A_IWL<1561> A_IWL<1560> A_IWL<1559> A_IWL<1558> A_IWL<1557> A_IWL<1556> A_IWL<1555> A_IWL<1554> A_IWL<1553> A_IWL<1552> A_IWL<1551> A_IWL<1550> A_IWL<1549> A_IWL<1548> A_IWL<1547> A_IWL<1546> A_IWL<1545> A_IWL<1544> A_IWL<1543> A_IWL<1542> A_IWL<1541> A_IWL<1540> A_IWL<1539> A_IWL<1538> A_IWL<1537> A_IWL<1536> A_IWL<2047> A_IWL<2046> A_IWL<2045> A_IWL<2044> A_IWL<2043> A_IWL<2042> A_IWL<2041> A_IWL<2040> A_IWL<2039> A_IWL<2038> A_IWL<2037> A_IWL<2036> A_IWL<2035> A_IWL<2034> A_IWL<2033> A_IWL<2032> A_IWL<2031> A_IWL<2030> A_IWL<2029> A_IWL<2028> A_IWL<2027> A_IWL<2026> A_IWL<2025> A_IWL<2024> A_IWL<2023> A_IWL<2022> A_IWL<2021> A_IWL<2020> A_IWL<2019> A_IWL<2018> A_IWL<2017> A_IWL<2016> A_IWL<2015> A_IWL<2014> A_IWL<2013> A_IWL<2012> A_IWL<2011> A_IWL<2010> A_IWL<2009> A_IWL<2008> A_IWL<2007> A_IWL<2006> A_IWL<2005> A_IWL<2004> A_IWL<2003> A_IWL<2002> A_IWL<2001> A_IWL<2000> A_IWL<1999> A_IWL<1998> A_IWL<1997> A_IWL<1996> A_IWL<1995> A_IWL<1994> A_IWL<1993> A_IWL<1992> A_IWL<1991> A_IWL<1990> A_IWL<1989> A_IWL<1988> A_IWL<1987> A_IWL<1986> A_IWL<1985> A_IWL<1984> A_IWL<1983> A_IWL<1982> A_IWL<1981> A_IWL<1980> A_IWL<1979> A_IWL<1978> A_IWL<1977> A_IWL<1976> A_IWL<1975> A_IWL<1974> A_IWL<1973> A_IWL<1972> A_IWL<1971> A_IWL<1970> A_IWL<1969> A_IWL<1968> A_IWL<1967> A_IWL<1966> A_IWL<1965> A_IWL<1964> A_IWL<1963> A_IWL<1962> A_IWL<1961> A_IWL<1960> A_IWL<1959> A_IWL<1958> A_IWL<1957> A_IWL<1956> A_IWL<1955> A_IWL<1954> A_IWL<1953> A_IWL<1952> A_IWL<1951> A_IWL<1950> A_IWL<1949> A_IWL<1948> A_IWL<1947> A_IWL<1946> A_IWL<1945> A_IWL<1944> A_IWL<1943> A_IWL<1942> A_IWL<1941> A_IWL<1940> A_IWL<1939> A_IWL<1938> A_IWL<1937> A_IWL<1936> A_IWL<1935> A_IWL<1934> A_IWL<1933> A_IWL<1932> A_IWL<1931> A_IWL<1930> A_IWL<1929> A_IWL<1928> A_IWL<1927> A_IWL<1926> A_IWL<1925> A_IWL<1924> A_IWL<1923> A_IWL<1922> A_IWL<1921> A_IWL<1920> A_IWL<1919> A_IWL<1918> A_IWL<1917> A_IWL<1916> A_IWL<1915> A_IWL<1914> A_IWL<1913> A_IWL<1912> A_IWL<1911> A_IWL<1910> A_IWL<1909> A_IWL<1908> A_IWL<1907> A_IWL<1906> A_IWL<1905> A_IWL<1904> A_IWL<1903> A_IWL<1902> A_IWL<1901> A_IWL<1900> A_IWL<1899> A_IWL<1898> A_IWL<1897> A_IWL<1896> A_IWL<1895> A_IWL<1894> A_IWL<1893> A_IWL<1892> A_IWL<1891> A_IWL<1890> A_IWL<1889> A_IWL<1888> A_IWL<1887> A_IWL<1886> A_IWL<1885> A_IWL<1884> A_IWL<1883> A_IWL<1882> A_IWL<1881> A_IWL<1880> A_IWL<1879> A_IWL<1878> A_IWL<1877> A_IWL<1876> A_IWL<1875> A_IWL<1874> A_IWL<1873> A_IWL<1872> A_IWL<1871> A_IWL<1870> A_IWL<1869> A_IWL<1868> A_IWL<1867> A_IWL<1866> A_IWL<1865> A_IWL<1864> A_IWL<1863> A_IWL<1862> A_IWL<1861> A_IWL<1860> A_IWL<1859> A_IWL<1858> A_IWL<1857> A_IWL<1856> A_IWL<1855> A_IWL<1854> A_IWL<1853> A_IWL<1852> A_IWL<1851> A_IWL<1850> A_IWL<1849> A_IWL<1848> A_IWL<1847> A_IWL<1846> A_IWL<1845> A_IWL<1844> A_IWL<1843> A_IWL<1842> A_IWL<1841> A_IWL<1840> A_IWL<1839> A_IWL<1838> A_IWL<1837> A_IWL<1836> A_IWL<1835> A_IWL<1834> A_IWL<1833> A_IWL<1832> A_IWL<1831> A_IWL<1830> A_IWL<1829> A_IWL<1828> A_IWL<1827> A_IWL<1826> A_IWL<1825> A_IWL<1824> A_IWL<1823> A_IWL<1822> A_IWL<1821> A_IWL<1820> A_IWL<1819> A_IWL<1818> A_IWL<1817> A_IWL<1816> A_IWL<1815> A_IWL<1814> A_IWL<1813> A_IWL<1812> A_IWL<1811> A_IWL<1810> A_IWL<1809> A_IWL<1808> A_IWL<1807> A_IWL<1806> A_IWL<1805> A_IWL<1804> A_IWL<1803> A_IWL<1802> A_IWL<1801> A_IWL<1800> A_IWL<1799> A_IWL<1798> A_IWL<1797> A_IWL<1796> A_IWL<1795> A_IWL<1794> A_IWL<1793> A_IWL<1792> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<6> A_BLC<13> A_BLC<12> A_BLC_TOP<13> A_BLC_TOP<12> A_BLT<13> A_BLT<12> A_BLT_TOP<13> A_BLT_TOP<12> A_IWL<1535> A_IWL<1534> A_IWL<1533> A_IWL<1532> A_IWL<1531> A_IWL<1530> A_IWL<1529> A_IWL<1528> A_IWL<1527> A_IWL<1526> A_IWL<1525> A_IWL<1524> A_IWL<1523> A_IWL<1522> A_IWL<1521> A_IWL<1520> A_IWL<1519> A_IWL<1518> A_IWL<1517> A_IWL<1516> A_IWL<1515> A_IWL<1514> A_IWL<1513> A_IWL<1512> A_IWL<1511> A_IWL<1510> A_IWL<1509> A_IWL<1508> A_IWL<1507> A_IWL<1506> A_IWL<1505> A_IWL<1504> A_IWL<1503> A_IWL<1502> A_IWL<1501> A_IWL<1500> A_IWL<1499> A_IWL<1498> A_IWL<1497> A_IWL<1496> A_IWL<1495> A_IWL<1494> A_IWL<1493> A_IWL<1492> A_IWL<1491> A_IWL<1490> A_IWL<1489> A_IWL<1488> A_IWL<1487> A_IWL<1486> A_IWL<1485> A_IWL<1484> A_IWL<1483> A_IWL<1482> A_IWL<1481> A_IWL<1480> A_IWL<1479> A_IWL<1478> A_IWL<1477> A_IWL<1476> A_IWL<1475> A_IWL<1474> A_IWL<1473> A_IWL<1472> A_IWL<1471> A_IWL<1470> A_IWL<1469> A_IWL<1468> A_IWL<1467> A_IWL<1466> A_IWL<1465> A_IWL<1464> A_IWL<1463> A_IWL<1462> A_IWL<1461> A_IWL<1460> A_IWL<1459> A_IWL<1458> A_IWL<1457> A_IWL<1456> A_IWL<1455> A_IWL<1454> A_IWL<1453> A_IWL<1452> A_IWL<1451> A_IWL<1450> A_IWL<1449> A_IWL<1448> A_IWL<1447> A_IWL<1446> A_IWL<1445> A_IWL<1444> A_IWL<1443> A_IWL<1442> A_IWL<1441> A_IWL<1440> A_IWL<1439> A_IWL<1438> A_IWL<1437> A_IWL<1436> A_IWL<1435> A_IWL<1434> A_IWL<1433> A_IWL<1432> A_IWL<1431> A_IWL<1430> A_IWL<1429> A_IWL<1428> A_IWL<1427> A_IWL<1426> A_IWL<1425> A_IWL<1424> A_IWL<1423> A_IWL<1422> A_IWL<1421> A_IWL<1420> A_IWL<1419> A_IWL<1418> A_IWL<1417> A_IWL<1416> A_IWL<1415> A_IWL<1414> A_IWL<1413> A_IWL<1412> A_IWL<1411> A_IWL<1410> A_IWL<1409> A_IWL<1408> A_IWL<1407> A_IWL<1406> A_IWL<1405> A_IWL<1404> A_IWL<1403> A_IWL<1402> A_IWL<1401> A_IWL<1400> A_IWL<1399> A_IWL<1398> A_IWL<1397> A_IWL<1396> A_IWL<1395> A_IWL<1394> A_IWL<1393> A_IWL<1392> A_IWL<1391> A_IWL<1390> A_IWL<1389> A_IWL<1388> A_IWL<1387> A_IWL<1386> A_IWL<1385> A_IWL<1384> A_IWL<1383> A_IWL<1382> A_IWL<1381> A_IWL<1380> A_IWL<1379> A_IWL<1378> A_IWL<1377> A_IWL<1376> A_IWL<1375> A_IWL<1374> A_IWL<1373> A_IWL<1372> A_IWL<1371> A_IWL<1370> A_IWL<1369> A_IWL<1368> A_IWL<1367> A_IWL<1366> A_IWL<1365> A_IWL<1364> A_IWL<1363> A_IWL<1362> A_IWL<1361> A_IWL<1360> A_IWL<1359> A_IWL<1358> A_IWL<1357> A_IWL<1356> A_IWL<1355> A_IWL<1354> A_IWL<1353> A_IWL<1352> A_IWL<1351> A_IWL<1350> A_IWL<1349> A_IWL<1348> A_IWL<1347> A_IWL<1346> A_IWL<1345> A_IWL<1344> A_IWL<1343> A_IWL<1342> A_IWL<1341> A_IWL<1340> A_IWL<1339> A_IWL<1338> A_IWL<1337> A_IWL<1336> A_IWL<1335> A_IWL<1334> A_IWL<1333> A_IWL<1332> A_IWL<1331> A_IWL<1330> A_IWL<1329> A_IWL<1328> A_IWL<1327> A_IWL<1326> A_IWL<1325> A_IWL<1324> A_IWL<1323> A_IWL<1322> A_IWL<1321> A_IWL<1320> A_IWL<1319> A_IWL<1318> A_IWL<1317> A_IWL<1316> A_IWL<1315> A_IWL<1314> A_IWL<1313> A_IWL<1312> A_IWL<1311> A_IWL<1310> A_IWL<1309> A_IWL<1308> A_IWL<1307> A_IWL<1306> A_IWL<1305> A_IWL<1304> A_IWL<1303> A_IWL<1302> A_IWL<1301> A_IWL<1300> A_IWL<1299> A_IWL<1298> A_IWL<1297> A_IWL<1296> A_IWL<1295> A_IWL<1294> A_IWL<1293> A_IWL<1292> A_IWL<1291> A_IWL<1290> A_IWL<1289> A_IWL<1288> A_IWL<1287> A_IWL<1286> A_IWL<1285> A_IWL<1284> A_IWL<1283> A_IWL<1282> A_IWL<1281> A_IWL<1280> A_IWL<1791> A_IWL<1790> A_IWL<1789> A_IWL<1788> A_IWL<1787> A_IWL<1786> A_IWL<1785> A_IWL<1784> A_IWL<1783> A_IWL<1782> A_IWL<1781> A_IWL<1780> A_IWL<1779> A_IWL<1778> A_IWL<1777> A_IWL<1776> A_IWL<1775> A_IWL<1774> A_IWL<1773> A_IWL<1772> A_IWL<1771> A_IWL<1770> A_IWL<1769> A_IWL<1768> A_IWL<1767> A_IWL<1766> A_IWL<1765> A_IWL<1764> A_IWL<1763> A_IWL<1762> A_IWL<1761> A_IWL<1760> A_IWL<1759> A_IWL<1758> A_IWL<1757> A_IWL<1756> A_IWL<1755> A_IWL<1754> A_IWL<1753> A_IWL<1752> A_IWL<1751> A_IWL<1750> A_IWL<1749> A_IWL<1748> A_IWL<1747> A_IWL<1746> A_IWL<1745> A_IWL<1744> A_IWL<1743> A_IWL<1742> A_IWL<1741> A_IWL<1740> A_IWL<1739> A_IWL<1738> A_IWL<1737> A_IWL<1736> A_IWL<1735> A_IWL<1734> A_IWL<1733> A_IWL<1732> A_IWL<1731> A_IWL<1730> A_IWL<1729> A_IWL<1728> A_IWL<1727> A_IWL<1726> A_IWL<1725> A_IWL<1724> A_IWL<1723> A_IWL<1722> A_IWL<1721> A_IWL<1720> A_IWL<1719> A_IWL<1718> A_IWL<1717> A_IWL<1716> A_IWL<1715> A_IWL<1714> A_IWL<1713> A_IWL<1712> A_IWL<1711> A_IWL<1710> A_IWL<1709> A_IWL<1708> A_IWL<1707> A_IWL<1706> A_IWL<1705> A_IWL<1704> A_IWL<1703> A_IWL<1702> A_IWL<1701> A_IWL<1700> A_IWL<1699> A_IWL<1698> A_IWL<1697> A_IWL<1696> A_IWL<1695> A_IWL<1694> A_IWL<1693> A_IWL<1692> A_IWL<1691> A_IWL<1690> A_IWL<1689> A_IWL<1688> A_IWL<1687> A_IWL<1686> A_IWL<1685> A_IWL<1684> A_IWL<1683> A_IWL<1682> A_IWL<1681> A_IWL<1680> A_IWL<1679> A_IWL<1678> A_IWL<1677> A_IWL<1676> A_IWL<1675> A_IWL<1674> A_IWL<1673> A_IWL<1672> A_IWL<1671> A_IWL<1670> A_IWL<1669> A_IWL<1668> A_IWL<1667> A_IWL<1666> A_IWL<1665> A_IWL<1664> A_IWL<1663> A_IWL<1662> A_IWL<1661> A_IWL<1660> A_IWL<1659> A_IWL<1658> A_IWL<1657> A_IWL<1656> A_IWL<1655> A_IWL<1654> A_IWL<1653> A_IWL<1652> A_IWL<1651> A_IWL<1650> A_IWL<1649> A_IWL<1648> A_IWL<1647> A_IWL<1646> A_IWL<1645> A_IWL<1644> A_IWL<1643> A_IWL<1642> A_IWL<1641> A_IWL<1640> A_IWL<1639> A_IWL<1638> A_IWL<1637> A_IWL<1636> A_IWL<1635> A_IWL<1634> A_IWL<1633> A_IWL<1632> A_IWL<1631> A_IWL<1630> A_IWL<1629> A_IWL<1628> A_IWL<1627> A_IWL<1626> A_IWL<1625> A_IWL<1624> A_IWL<1623> A_IWL<1622> A_IWL<1621> A_IWL<1620> A_IWL<1619> A_IWL<1618> A_IWL<1617> A_IWL<1616> A_IWL<1615> A_IWL<1614> A_IWL<1613> A_IWL<1612> A_IWL<1611> A_IWL<1610> A_IWL<1609> A_IWL<1608> A_IWL<1607> A_IWL<1606> A_IWL<1605> A_IWL<1604> A_IWL<1603> A_IWL<1602> A_IWL<1601> A_IWL<1600> A_IWL<1599> A_IWL<1598> A_IWL<1597> A_IWL<1596> A_IWL<1595> A_IWL<1594> A_IWL<1593> A_IWL<1592> A_IWL<1591> A_IWL<1590> A_IWL<1589> A_IWL<1588> A_IWL<1587> A_IWL<1586> A_IWL<1585> A_IWL<1584> A_IWL<1583> A_IWL<1582> A_IWL<1581> A_IWL<1580> A_IWL<1579> A_IWL<1578> A_IWL<1577> A_IWL<1576> A_IWL<1575> A_IWL<1574> A_IWL<1573> A_IWL<1572> A_IWL<1571> A_IWL<1570> A_IWL<1569> A_IWL<1568> A_IWL<1567> A_IWL<1566> A_IWL<1565> A_IWL<1564> A_IWL<1563> A_IWL<1562> A_IWL<1561> A_IWL<1560> A_IWL<1559> A_IWL<1558> A_IWL<1557> A_IWL<1556> A_IWL<1555> A_IWL<1554> A_IWL<1553> A_IWL<1552> A_IWL<1551> A_IWL<1550> A_IWL<1549> A_IWL<1548> A_IWL<1547> A_IWL<1546> A_IWL<1545> A_IWL<1544> A_IWL<1543> A_IWL<1542> A_IWL<1541> A_IWL<1540> A_IWL<1539> A_IWL<1538> A_IWL<1537> A_IWL<1536> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<5> A_BLC<11> A_BLC<10> A_BLC_TOP<11> A_BLC_TOP<10> A_BLT<11> A_BLT<10> A_BLT_TOP<11> A_BLT_TOP<10> A_IWL<1279> A_IWL<1278> A_IWL<1277> A_IWL<1276> A_IWL<1275> A_IWL<1274> A_IWL<1273> A_IWL<1272> A_IWL<1271> A_IWL<1270> A_IWL<1269> A_IWL<1268> A_IWL<1267> A_IWL<1266> A_IWL<1265> A_IWL<1264> A_IWL<1263> A_IWL<1262> A_IWL<1261> A_IWL<1260> A_IWL<1259> A_IWL<1258> A_IWL<1257> A_IWL<1256> A_IWL<1255> A_IWL<1254> A_IWL<1253> A_IWL<1252> A_IWL<1251> A_IWL<1250> A_IWL<1249> A_IWL<1248> A_IWL<1247> A_IWL<1246> A_IWL<1245> A_IWL<1244> A_IWL<1243> A_IWL<1242> A_IWL<1241> A_IWL<1240> A_IWL<1239> A_IWL<1238> A_IWL<1237> A_IWL<1236> A_IWL<1235> A_IWL<1234> A_IWL<1233> A_IWL<1232> A_IWL<1231> A_IWL<1230> A_IWL<1229> A_IWL<1228> A_IWL<1227> A_IWL<1226> A_IWL<1225> A_IWL<1224> A_IWL<1223> A_IWL<1222> A_IWL<1221> A_IWL<1220> A_IWL<1219> A_IWL<1218> A_IWL<1217> A_IWL<1216> A_IWL<1215> A_IWL<1214> A_IWL<1213> A_IWL<1212> A_IWL<1211> A_IWL<1210> A_IWL<1209> A_IWL<1208> A_IWL<1207> A_IWL<1206> A_IWL<1205> A_IWL<1204> A_IWL<1203> A_IWL<1202> A_IWL<1201> A_IWL<1200> A_IWL<1199> A_IWL<1198> A_IWL<1197> A_IWL<1196> A_IWL<1195> A_IWL<1194> A_IWL<1193> A_IWL<1192> A_IWL<1191> A_IWL<1190> A_IWL<1189> A_IWL<1188> A_IWL<1187> A_IWL<1186> A_IWL<1185> A_IWL<1184> A_IWL<1183> A_IWL<1182> A_IWL<1181> A_IWL<1180> A_IWL<1179> A_IWL<1178> A_IWL<1177> A_IWL<1176> A_IWL<1175> A_IWL<1174> A_IWL<1173> A_IWL<1172> A_IWL<1171> A_IWL<1170> A_IWL<1169> A_IWL<1168> A_IWL<1167> A_IWL<1166> A_IWL<1165> A_IWL<1164> A_IWL<1163> A_IWL<1162> A_IWL<1161> A_IWL<1160> A_IWL<1159> A_IWL<1158> A_IWL<1157> A_IWL<1156> A_IWL<1155> A_IWL<1154> A_IWL<1153> A_IWL<1152> A_IWL<1151> A_IWL<1150> A_IWL<1149> A_IWL<1148> A_IWL<1147> A_IWL<1146> A_IWL<1145> A_IWL<1144> A_IWL<1143> A_IWL<1142> A_IWL<1141> A_IWL<1140> A_IWL<1139> A_IWL<1138> A_IWL<1137> A_IWL<1136> A_IWL<1135> A_IWL<1134> A_IWL<1133> A_IWL<1132> A_IWL<1131> A_IWL<1130> A_IWL<1129> A_IWL<1128> A_IWL<1127> A_IWL<1126> A_IWL<1125> A_IWL<1124> A_IWL<1123> A_IWL<1122> A_IWL<1121> A_IWL<1120> A_IWL<1119> A_IWL<1118> A_IWL<1117> A_IWL<1116> A_IWL<1115> A_IWL<1114> A_IWL<1113> A_IWL<1112> A_IWL<1111> A_IWL<1110> A_IWL<1109> A_IWL<1108> A_IWL<1107> A_IWL<1106> A_IWL<1105> A_IWL<1104> A_IWL<1103> A_IWL<1102> A_IWL<1101> A_IWL<1100> A_IWL<1099> A_IWL<1098> A_IWL<1097> A_IWL<1096> A_IWL<1095> A_IWL<1094> A_IWL<1093> A_IWL<1092> A_IWL<1091> A_IWL<1090> A_IWL<1089> A_IWL<1088> A_IWL<1087> A_IWL<1086> A_IWL<1085> A_IWL<1084> A_IWL<1083> A_IWL<1082> A_IWL<1081> A_IWL<1080> A_IWL<1079> A_IWL<1078> A_IWL<1077> A_IWL<1076> A_IWL<1075> A_IWL<1074> A_IWL<1073> A_IWL<1072> A_IWL<1071> A_IWL<1070> A_IWL<1069> A_IWL<1068> A_IWL<1067> A_IWL<1066> A_IWL<1065> A_IWL<1064> A_IWL<1063> A_IWL<1062> A_IWL<1061> A_IWL<1060> A_IWL<1059> A_IWL<1058> A_IWL<1057> A_IWL<1056> A_IWL<1055> A_IWL<1054> A_IWL<1053> A_IWL<1052> A_IWL<1051> A_IWL<1050> A_IWL<1049> A_IWL<1048> A_IWL<1047> A_IWL<1046> A_IWL<1045> A_IWL<1044> A_IWL<1043> A_IWL<1042> A_IWL<1041> A_IWL<1040> A_IWL<1039> A_IWL<1038> A_IWL<1037> A_IWL<1036> A_IWL<1035> A_IWL<1034> A_IWL<1033> A_IWL<1032> A_IWL<1031> A_IWL<1030> A_IWL<1029> A_IWL<1028> A_IWL<1027> A_IWL<1026> A_IWL<1025> A_IWL<1024> A_IWL<1535> A_IWL<1534> A_IWL<1533> A_IWL<1532> A_IWL<1531> A_IWL<1530> A_IWL<1529> A_IWL<1528> A_IWL<1527> A_IWL<1526> A_IWL<1525> A_IWL<1524> A_IWL<1523> A_IWL<1522> A_IWL<1521> A_IWL<1520> A_IWL<1519> A_IWL<1518> A_IWL<1517> A_IWL<1516> A_IWL<1515> A_IWL<1514> A_IWL<1513> A_IWL<1512> A_IWL<1511> A_IWL<1510> A_IWL<1509> A_IWL<1508> A_IWL<1507> A_IWL<1506> A_IWL<1505> A_IWL<1504> A_IWL<1503> A_IWL<1502> A_IWL<1501> A_IWL<1500> A_IWL<1499> A_IWL<1498> A_IWL<1497> A_IWL<1496> A_IWL<1495> A_IWL<1494> A_IWL<1493> A_IWL<1492> A_IWL<1491> A_IWL<1490> A_IWL<1489> A_IWL<1488> A_IWL<1487> A_IWL<1486> A_IWL<1485> A_IWL<1484> A_IWL<1483> A_IWL<1482> A_IWL<1481> A_IWL<1480> A_IWL<1479> A_IWL<1478> A_IWL<1477> A_IWL<1476> A_IWL<1475> A_IWL<1474> A_IWL<1473> A_IWL<1472> A_IWL<1471> A_IWL<1470> A_IWL<1469> A_IWL<1468> A_IWL<1467> A_IWL<1466> A_IWL<1465> A_IWL<1464> A_IWL<1463> A_IWL<1462> A_IWL<1461> A_IWL<1460> A_IWL<1459> A_IWL<1458> A_IWL<1457> A_IWL<1456> A_IWL<1455> A_IWL<1454> A_IWL<1453> A_IWL<1452> A_IWL<1451> A_IWL<1450> A_IWL<1449> A_IWL<1448> A_IWL<1447> A_IWL<1446> A_IWL<1445> A_IWL<1444> A_IWL<1443> A_IWL<1442> A_IWL<1441> A_IWL<1440> A_IWL<1439> A_IWL<1438> A_IWL<1437> A_IWL<1436> A_IWL<1435> A_IWL<1434> A_IWL<1433> A_IWL<1432> A_IWL<1431> A_IWL<1430> A_IWL<1429> A_IWL<1428> A_IWL<1427> A_IWL<1426> A_IWL<1425> A_IWL<1424> A_IWL<1423> A_IWL<1422> A_IWL<1421> A_IWL<1420> A_IWL<1419> A_IWL<1418> A_IWL<1417> A_IWL<1416> A_IWL<1415> A_IWL<1414> A_IWL<1413> A_IWL<1412> A_IWL<1411> A_IWL<1410> A_IWL<1409> A_IWL<1408> A_IWL<1407> A_IWL<1406> A_IWL<1405> A_IWL<1404> A_IWL<1403> A_IWL<1402> A_IWL<1401> A_IWL<1400> A_IWL<1399> A_IWL<1398> A_IWL<1397> A_IWL<1396> A_IWL<1395> A_IWL<1394> A_IWL<1393> A_IWL<1392> A_IWL<1391> A_IWL<1390> A_IWL<1389> A_IWL<1388> A_IWL<1387> A_IWL<1386> A_IWL<1385> A_IWL<1384> A_IWL<1383> A_IWL<1382> A_IWL<1381> A_IWL<1380> A_IWL<1379> A_IWL<1378> A_IWL<1377> A_IWL<1376> A_IWL<1375> A_IWL<1374> A_IWL<1373> A_IWL<1372> A_IWL<1371> A_IWL<1370> A_IWL<1369> A_IWL<1368> A_IWL<1367> A_IWL<1366> A_IWL<1365> A_IWL<1364> A_IWL<1363> A_IWL<1362> A_IWL<1361> A_IWL<1360> A_IWL<1359> A_IWL<1358> A_IWL<1357> A_IWL<1356> A_IWL<1355> A_IWL<1354> A_IWL<1353> A_IWL<1352> A_IWL<1351> A_IWL<1350> A_IWL<1349> A_IWL<1348> A_IWL<1347> A_IWL<1346> A_IWL<1345> A_IWL<1344> A_IWL<1343> A_IWL<1342> A_IWL<1341> A_IWL<1340> A_IWL<1339> A_IWL<1338> A_IWL<1337> A_IWL<1336> A_IWL<1335> A_IWL<1334> A_IWL<1333> A_IWL<1332> A_IWL<1331> A_IWL<1330> A_IWL<1329> A_IWL<1328> A_IWL<1327> A_IWL<1326> A_IWL<1325> A_IWL<1324> A_IWL<1323> A_IWL<1322> A_IWL<1321> A_IWL<1320> A_IWL<1319> A_IWL<1318> A_IWL<1317> A_IWL<1316> A_IWL<1315> A_IWL<1314> A_IWL<1313> A_IWL<1312> A_IWL<1311> A_IWL<1310> A_IWL<1309> A_IWL<1308> A_IWL<1307> A_IWL<1306> A_IWL<1305> A_IWL<1304> A_IWL<1303> A_IWL<1302> A_IWL<1301> A_IWL<1300> A_IWL<1299> A_IWL<1298> A_IWL<1297> A_IWL<1296> A_IWL<1295> A_IWL<1294> A_IWL<1293> A_IWL<1292> A_IWL<1291> A_IWL<1290> A_IWL<1289> A_IWL<1288> A_IWL<1287> A_IWL<1286> A_IWL<1285> A_IWL<1284> A_IWL<1283> A_IWL<1282> A_IWL<1281> A_IWL<1280> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<4> A_BLC<9> A_BLC<8> A_BLC_TOP<9> A_BLC_TOP<8> A_BLT<9> A_BLT<8> A_BLT_TOP<9> A_BLT_TOP<8> A_IWL<1023> A_IWL<1022> A_IWL<1021> A_IWL<1020> A_IWL<1019> A_IWL<1018> A_IWL<1017> A_IWL<1016> A_IWL<1015> A_IWL<1014> A_IWL<1013> A_IWL<1012> A_IWL<1011> A_IWL<1010> A_IWL<1009> A_IWL<1008> A_IWL<1007> A_IWL<1006> A_IWL<1005> A_IWL<1004> A_IWL<1003> A_IWL<1002> A_IWL<1001> A_IWL<1000> A_IWL<999> A_IWL<998> A_IWL<997> A_IWL<996> A_IWL<995> A_IWL<994> A_IWL<993> A_IWL<992> A_IWL<991> A_IWL<990> A_IWL<989> A_IWL<988> A_IWL<987> A_IWL<986> A_IWL<985> A_IWL<984> A_IWL<983> A_IWL<982> A_IWL<981> A_IWL<980> A_IWL<979> A_IWL<978> A_IWL<977> A_IWL<976> A_IWL<975> A_IWL<974> A_IWL<973> A_IWL<972> A_IWL<971> A_IWL<970> A_IWL<969> A_IWL<968> A_IWL<967> A_IWL<966> A_IWL<965> A_IWL<964> A_IWL<963> A_IWL<962> A_IWL<961> A_IWL<960> A_IWL<959> A_IWL<958> A_IWL<957> A_IWL<956> A_IWL<955> A_IWL<954> A_IWL<953> A_IWL<952> A_IWL<951> A_IWL<950> A_IWL<949> A_IWL<948> A_IWL<947> A_IWL<946> A_IWL<945> A_IWL<944> A_IWL<943> A_IWL<942> A_IWL<941> A_IWL<940> A_IWL<939> A_IWL<938> A_IWL<937> A_IWL<936> A_IWL<935> A_IWL<934> A_IWL<933> A_IWL<932> A_IWL<931> A_IWL<930> A_IWL<929> A_IWL<928> A_IWL<927> A_IWL<926> A_IWL<925> A_IWL<924> A_IWL<923> A_IWL<922> A_IWL<921> A_IWL<920> A_IWL<919> A_IWL<918> A_IWL<917> A_IWL<916> A_IWL<915> A_IWL<914> A_IWL<913> A_IWL<912> A_IWL<911> A_IWL<910> A_IWL<909> A_IWL<908> A_IWL<907> A_IWL<906> A_IWL<905> A_IWL<904> A_IWL<903> A_IWL<902> A_IWL<901> A_IWL<900> A_IWL<899> A_IWL<898> A_IWL<897> A_IWL<896> A_IWL<895> A_IWL<894> A_IWL<893> A_IWL<892> A_IWL<891> A_IWL<890> A_IWL<889> A_IWL<888> A_IWL<887> A_IWL<886> A_IWL<885> A_IWL<884> A_IWL<883> A_IWL<882> A_IWL<881> A_IWL<880> A_IWL<879> A_IWL<878> A_IWL<877> A_IWL<876> A_IWL<875> A_IWL<874> A_IWL<873> A_IWL<872> A_IWL<871> A_IWL<870> A_IWL<869> A_IWL<868> A_IWL<867> A_IWL<866> A_IWL<865> A_IWL<864> A_IWL<863> A_IWL<862> A_IWL<861> A_IWL<860> A_IWL<859> A_IWL<858> A_IWL<857> A_IWL<856> A_IWL<855> A_IWL<854> A_IWL<853> A_IWL<852> A_IWL<851> A_IWL<850> A_IWL<849> A_IWL<848> A_IWL<847> A_IWL<846> A_IWL<845> A_IWL<844> A_IWL<843> A_IWL<842> A_IWL<841> A_IWL<840> A_IWL<839> A_IWL<838> A_IWL<837> A_IWL<836> A_IWL<835> A_IWL<834> A_IWL<833> A_IWL<832> A_IWL<831> A_IWL<830> A_IWL<829> A_IWL<828> A_IWL<827> A_IWL<826> A_IWL<825> A_IWL<824> A_IWL<823> A_IWL<822> A_IWL<821> A_IWL<820> A_IWL<819> A_IWL<818> A_IWL<817> A_IWL<816> A_IWL<815> A_IWL<814> A_IWL<813> A_IWL<812> A_IWL<811> A_IWL<810> A_IWL<809> A_IWL<808> A_IWL<807> A_IWL<806> A_IWL<805> A_IWL<804> A_IWL<803> A_IWL<802> A_IWL<801> A_IWL<800> A_IWL<799> A_IWL<798> A_IWL<797> A_IWL<796> A_IWL<795> A_IWL<794> A_IWL<793> A_IWL<792> A_IWL<791> A_IWL<790> A_IWL<789> A_IWL<788> A_IWL<787> A_IWL<786> A_IWL<785> A_IWL<784> A_IWL<783> A_IWL<782> A_IWL<781> A_IWL<780> A_IWL<779> A_IWL<778> A_IWL<777> A_IWL<776> A_IWL<775> A_IWL<774> A_IWL<773> A_IWL<772> A_IWL<771> A_IWL<770> A_IWL<769> A_IWL<768> A_IWL<1279> A_IWL<1278> A_IWL<1277> A_IWL<1276> A_IWL<1275> A_IWL<1274> A_IWL<1273> A_IWL<1272> A_IWL<1271> A_IWL<1270> A_IWL<1269> A_IWL<1268> A_IWL<1267> A_IWL<1266> A_IWL<1265> A_IWL<1264> A_IWL<1263> A_IWL<1262> A_IWL<1261> A_IWL<1260> A_IWL<1259> A_IWL<1258> A_IWL<1257> A_IWL<1256> A_IWL<1255> A_IWL<1254> A_IWL<1253> A_IWL<1252> A_IWL<1251> A_IWL<1250> A_IWL<1249> A_IWL<1248> A_IWL<1247> A_IWL<1246> A_IWL<1245> A_IWL<1244> A_IWL<1243> A_IWL<1242> A_IWL<1241> A_IWL<1240> A_IWL<1239> A_IWL<1238> A_IWL<1237> A_IWL<1236> A_IWL<1235> A_IWL<1234> A_IWL<1233> A_IWL<1232> A_IWL<1231> A_IWL<1230> A_IWL<1229> A_IWL<1228> A_IWL<1227> A_IWL<1226> A_IWL<1225> A_IWL<1224> A_IWL<1223> A_IWL<1222> A_IWL<1221> A_IWL<1220> A_IWL<1219> A_IWL<1218> A_IWL<1217> A_IWL<1216> A_IWL<1215> A_IWL<1214> A_IWL<1213> A_IWL<1212> A_IWL<1211> A_IWL<1210> A_IWL<1209> A_IWL<1208> A_IWL<1207> A_IWL<1206> A_IWL<1205> A_IWL<1204> A_IWL<1203> A_IWL<1202> A_IWL<1201> A_IWL<1200> A_IWL<1199> A_IWL<1198> A_IWL<1197> A_IWL<1196> A_IWL<1195> A_IWL<1194> A_IWL<1193> A_IWL<1192> A_IWL<1191> A_IWL<1190> A_IWL<1189> A_IWL<1188> A_IWL<1187> A_IWL<1186> A_IWL<1185> A_IWL<1184> A_IWL<1183> A_IWL<1182> A_IWL<1181> A_IWL<1180> A_IWL<1179> A_IWL<1178> A_IWL<1177> A_IWL<1176> A_IWL<1175> A_IWL<1174> A_IWL<1173> A_IWL<1172> A_IWL<1171> A_IWL<1170> A_IWL<1169> A_IWL<1168> A_IWL<1167> A_IWL<1166> A_IWL<1165> A_IWL<1164> A_IWL<1163> A_IWL<1162> A_IWL<1161> A_IWL<1160> A_IWL<1159> A_IWL<1158> A_IWL<1157> A_IWL<1156> A_IWL<1155> A_IWL<1154> A_IWL<1153> A_IWL<1152> A_IWL<1151> A_IWL<1150> A_IWL<1149> A_IWL<1148> A_IWL<1147> A_IWL<1146> A_IWL<1145> A_IWL<1144> A_IWL<1143> A_IWL<1142> A_IWL<1141> A_IWL<1140> A_IWL<1139> A_IWL<1138> A_IWL<1137> A_IWL<1136> A_IWL<1135> A_IWL<1134> A_IWL<1133> A_IWL<1132> A_IWL<1131> A_IWL<1130> A_IWL<1129> A_IWL<1128> A_IWL<1127> A_IWL<1126> A_IWL<1125> A_IWL<1124> A_IWL<1123> A_IWL<1122> A_IWL<1121> A_IWL<1120> A_IWL<1119> A_IWL<1118> A_IWL<1117> A_IWL<1116> A_IWL<1115> A_IWL<1114> A_IWL<1113> A_IWL<1112> A_IWL<1111> A_IWL<1110> A_IWL<1109> A_IWL<1108> A_IWL<1107> A_IWL<1106> A_IWL<1105> A_IWL<1104> A_IWL<1103> A_IWL<1102> A_IWL<1101> A_IWL<1100> A_IWL<1099> A_IWL<1098> A_IWL<1097> A_IWL<1096> A_IWL<1095> A_IWL<1094> A_IWL<1093> A_IWL<1092> A_IWL<1091> A_IWL<1090> A_IWL<1089> A_IWL<1088> A_IWL<1087> A_IWL<1086> A_IWL<1085> A_IWL<1084> A_IWL<1083> A_IWL<1082> A_IWL<1081> A_IWL<1080> A_IWL<1079> A_IWL<1078> A_IWL<1077> A_IWL<1076> A_IWL<1075> A_IWL<1074> A_IWL<1073> A_IWL<1072> A_IWL<1071> A_IWL<1070> A_IWL<1069> A_IWL<1068> A_IWL<1067> A_IWL<1066> A_IWL<1065> A_IWL<1064> A_IWL<1063> A_IWL<1062> A_IWL<1061> A_IWL<1060> A_IWL<1059> A_IWL<1058> A_IWL<1057> A_IWL<1056> A_IWL<1055> A_IWL<1054> A_IWL<1053> A_IWL<1052> A_IWL<1051> A_IWL<1050> A_IWL<1049> A_IWL<1048> A_IWL<1047> A_IWL<1046> A_IWL<1045> A_IWL<1044> A_IWL<1043> A_IWL<1042> A_IWL<1041> A_IWL<1040> A_IWL<1039> A_IWL<1038> A_IWL<1037> A_IWL<1036> A_IWL<1035> A_IWL<1034> A_IWL<1033> A_IWL<1032> A_IWL<1031> A_IWL<1030> A_IWL<1029> A_IWL<1028> A_IWL<1027> A_IWL<1026> A_IWL<1025> A_IWL<1024> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<3> A_BLC<7> A_BLC<6> A_BLC_TOP<7> A_BLC_TOP<6> A_BLT<7> A_BLT<6> A_BLT_TOP<7> A_BLT_TOP<6> A_IWL<767> A_IWL<766> A_IWL<765> A_IWL<764> A_IWL<763> A_IWL<762> A_IWL<761> A_IWL<760> A_IWL<759> A_IWL<758> A_IWL<757> A_IWL<756> A_IWL<755> A_IWL<754> A_IWL<753> A_IWL<752> A_IWL<751> A_IWL<750> A_IWL<749> A_IWL<748> A_IWL<747> A_IWL<746> A_IWL<745> A_IWL<744> A_IWL<743> A_IWL<742> A_IWL<741> A_IWL<740> A_IWL<739> A_IWL<738> A_IWL<737> A_IWL<736> A_IWL<735> A_IWL<734> A_IWL<733> A_IWL<732> A_IWL<731> A_IWL<730> A_IWL<729> A_IWL<728> A_IWL<727> A_IWL<726> A_IWL<725> A_IWL<724> A_IWL<723> A_IWL<722> A_IWL<721> A_IWL<720> A_IWL<719> A_IWL<718> A_IWL<717> A_IWL<716> A_IWL<715> A_IWL<714> A_IWL<713> A_IWL<712> A_IWL<711> A_IWL<710> A_IWL<709> A_IWL<708> A_IWL<707> A_IWL<706> A_IWL<705> A_IWL<704> A_IWL<703> A_IWL<702> A_IWL<701> A_IWL<700> A_IWL<699> A_IWL<698> A_IWL<697> A_IWL<696> A_IWL<695> A_IWL<694> A_IWL<693> A_IWL<692> A_IWL<691> A_IWL<690> A_IWL<689> A_IWL<688> A_IWL<687> A_IWL<686> A_IWL<685> A_IWL<684> A_IWL<683> A_IWL<682> A_IWL<681> A_IWL<680> A_IWL<679> A_IWL<678> A_IWL<677> A_IWL<676> A_IWL<675> A_IWL<674> A_IWL<673> A_IWL<672> A_IWL<671> A_IWL<670> A_IWL<669> A_IWL<668> A_IWL<667> A_IWL<666> A_IWL<665> A_IWL<664> A_IWL<663> A_IWL<662> A_IWL<661> A_IWL<660> A_IWL<659> A_IWL<658> A_IWL<657> A_IWL<656> A_IWL<655> A_IWL<654> A_IWL<653> A_IWL<652> A_IWL<651> A_IWL<650> A_IWL<649> A_IWL<648> A_IWL<647> A_IWL<646> A_IWL<645> A_IWL<644> A_IWL<643> A_IWL<642> A_IWL<641> A_IWL<640> A_IWL<639> A_IWL<638> A_IWL<637> A_IWL<636> A_IWL<635> A_IWL<634> A_IWL<633> A_IWL<632> A_IWL<631> A_IWL<630> A_IWL<629> A_IWL<628> A_IWL<627> A_IWL<626> A_IWL<625> A_IWL<624> A_IWL<623> A_IWL<622> A_IWL<621> A_IWL<620> A_IWL<619> A_IWL<618> A_IWL<617> A_IWL<616> A_IWL<615> A_IWL<614> A_IWL<613> A_IWL<612> A_IWL<611> A_IWL<610> A_IWL<609> A_IWL<608> A_IWL<607> A_IWL<606> A_IWL<605> A_IWL<604> A_IWL<603> A_IWL<602> A_IWL<601> A_IWL<600> A_IWL<599> A_IWL<598> A_IWL<597> A_IWL<596> A_IWL<595> A_IWL<594> A_IWL<593> A_IWL<592> A_IWL<591> A_IWL<590> A_IWL<589> A_IWL<588> A_IWL<587> A_IWL<586> A_IWL<585> A_IWL<584> A_IWL<583> A_IWL<582> A_IWL<581> A_IWL<580> A_IWL<579> A_IWL<578> A_IWL<577> A_IWL<576> A_IWL<575> A_IWL<574> A_IWL<573> A_IWL<572> A_IWL<571> A_IWL<570> A_IWL<569> A_IWL<568> A_IWL<567> A_IWL<566> A_IWL<565> A_IWL<564> A_IWL<563> A_IWL<562> A_IWL<561> A_IWL<560> A_IWL<559> A_IWL<558> A_IWL<557> A_IWL<556> A_IWL<555> A_IWL<554> A_IWL<553> A_IWL<552> A_IWL<551> A_IWL<550> A_IWL<549> A_IWL<548> A_IWL<547> A_IWL<546> A_IWL<545> A_IWL<544> A_IWL<543> A_IWL<542> A_IWL<541> A_IWL<540> A_IWL<539> A_IWL<538> A_IWL<537> A_IWL<536> A_IWL<535> A_IWL<534> A_IWL<533> A_IWL<532> A_IWL<531> A_IWL<530> A_IWL<529> A_IWL<528> A_IWL<527> A_IWL<526> A_IWL<525> A_IWL<524> A_IWL<523> A_IWL<522> A_IWL<521> A_IWL<520> A_IWL<519> A_IWL<518> A_IWL<517> A_IWL<516> A_IWL<515> A_IWL<514> A_IWL<513> A_IWL<512> A_IWL<1023> A_IWL<1022> A_IWL<1021> A_IWL<1020> A_IWL<1019> A_IWL<1018> A_IWL<1017> A_IWL<1016> A_IWL<1015> A_IWL<1014> A_IWL<1013> A_IWL<1012> A_IWL<1011> A_IWL<1010> A_IWL<1009> A_IWL<1008> A_IWL<1007> A_IWL<1006> A_IWL<1005> A_IWL<1004> A_IWL<1003> A_IWL<1002> A_IWL<1001> A_IWL<1000> A_IWL<999> A_IWL<998> A_IWL<997> A_IWL<996> A_IWL<995> A_IWL<994> A_IWL<993> A_IWL<992> A_IWL<991> A_IWL<990> A_IWL<989> A_IWL<988> A_IWL<987> A_IWL<986> A_IWL<985> A_IWL<984> A_IWL<983> A_IWL<982> A_IWL<981> A_IWL<980> A_IWL<979> A_IWL<978> A_IWL<977> A_IWL<976> A_IWL<975> A_IWL<974> A_IWL<973> A_IWL<972> A_IWL<971> A_IWL<970> A_IWL<969> A_IWL<968> A_IWL<967> A_IWL<966> A_IWL<965> A_IWL<964> A_IWL<963> A_IWL<962> A_IWL<961> A_IWL<960> A_IWL<959> A_IWL<958> A_IWL<957> A_IWL<956> A_IWL<955> A_IWL<954> A_IWL<953> A_IWL<952> A_IWL<951> A_IWL<950> A_IWL<949> A_IWL<948> A_IWL<947> A_IWL<946> A_IWL<945> A_IWL<944> A_IWL<943> A_IWL<942> A_IWL<941> A_IWL<940> A_IWL<939> A_IWL<938> A_IWL<937> A_IWL<936> A_IWL<935> A_IWL<934> A_IWL<933> A_IWL<932> A_IWL<931> A_IWL<930> A_IWL<929> A_IWL<928> A_IWL<927> A_IWL<926> A_IWL<925> A_IWL<924> A_IWL<923> A_IWL<922> A_IWL<921> A_IWL<920> A_IWL<919> A_IWL<918> A_IWL<917> A_IWL<916> A_IWL<915> A_IWL<914> A_IWL<913> A_IWL<912> A_IWL<911> A_IWL<910> A_IWL<909> A_IWL<908> A_IWL<907> A_IWL<906> A_IWL<905> A_IWL<904> A_IWL<903> A_IWL<902> A_IWL<901> A_IWL<900> A_IWL<899> A_IWL<898> A_IWL<897> A_IWL<896> A_IWL<895> A_IWL<894> A_IWL<893> A_IWL<892> A_IWL<891> A_IWL<890> A_IWL<889> A_IWL<888> A_IWL<887> A_IWL<886> A_IWL<885> A_IWL<884> A_IWL<883> A_IWL<882> A_IWL<881> A_IWL<880> A_IWL<879> A_IWL<878> A_IWL<877> A_IWL<876> A_IWL<875> A_IWL<874> A_IWL<873> A_IWL<872> A_IWL<871> A_IWL<870> A_IWL<869> A_IWL<868> A_IWL<867> A_IWL<866> A_IWL<865> A_IWL<864> A_IWL<863> A_IWL<862> A_IWL<861> A_IWL<860> A_IWL<859> A_IWL<858> A_IWL<857> A_IWL<856> A_IWL<855> A_IWL<854> A_IWL<853> A_IWL<852> A_IWL<851> A_IWL<850> A_IWL<849> A_IWL<848> A_IWL<847> A_IWL<846> A_IWL<845> A_IWL<844> A_IWL<843> A_IWL<842> A_IWL<841> A_IWL<840> A_IWL<839> A_IWL<838> A_IWL<837> A_IWL<836> A_IWL<835> A_IWL<834> A_IWL<833> A_IWL<832> A_IWL<831> A_IWL<830> A_IWL<829> A_IWL<828> A_IWL<827> A_IWL<826> A_IWL<825> A_IWL<824> A_IWL<823> A_IWL<822> A_IWL<821> A_IWL<820> A_IWL<819> A_IWL<818> A_IWL<817> A_IWL<816> A_IWL<815> A_IWL<814> A_IWL<813> A_IWL<812> A_IWL<811> A_IWL<810> A_IWL<809> A_IWL<808> A_IWL<807> A_IWL<806> A_IWL<805> A_IWL<804> A_IWL<803> A_IWL<802> A_IWL<801> A_IWL<800> A_IWL<799> A_IWL<798> A_IWL<797> A_IWL<796> A_IWL<795> A_IWL<794> A_IWL<793> A_IWL<792> A_IWL<791> A_IWL<790> A_IWL<789> A_IWL<788> A_IWL<787> A_IWL<786> A_IWL<785> A_IWL<784> A_IWL<783> A_IWL<782> A_IWL<781> A_IWL<780> A_IWL<779> A_IWL<778> A_IWL<777> A_IWL<776> A_IWL<775> A_IWL<774> A_IWL<773> A_IWL<772> A_IWL<771> A_IWL<770> A_IWL<769> A_IWL<768> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<2> A_BLC<5> A_BLC<4> A_BLC_TOP<5> A_BLC_TOP<4> A_BLT<5> A_BLT<4> A_BLT_TOP<5> A_BLT_TOP<4> A_IWL<511> A_IWL<510> A_IWL<509> A_IWL<508> A_IWL<507> A_IWL<506> A_IWL<505> A_IWL<504> A_IWL<503> A_IWL<502> A_IWL<501> A_IWL<500> A_IWL<499> A_IWL<498> A_IWL<497> A_IWL<496> A_IWL<495> A_IWL<494> A_IWL<493> A_IWL<492> A_IWL<491> A_IWL<490> A_IWL<489> A_IWL<488> A_IWL<487> A_IWL<486> A_IWL<485> A_IWL<484> A_IWL<483> A_IWL<482> A_IWL<481> A_IWL<480> A_IWL<479> A_IWL<478> A_IWL<477> A_IWL<476> A_IWL<475> A_IWL<474> A_IWL<473> A_IWL<472> A_IWL<471> A_IWL<470> A_IWL<469> A_IWL<468> A_IWL<467> A_IWL<466> A_IWL<465> A_IWL<464> A_IWL<463> A_IWL<462> A_IWL<461> A_IWL<460> A_IWL<459> A_IWL<458> A_IWL<457> A_IWL<456> A_IWL<455> A_IWL<454> A_IWL<453> A_IWL<452> A_IWL<451> A_IWL<450> A_IWL<449> A_IWL<448> A_IWL<447> A_IWL<446> A_IWL<445> A_IWL<444> A_IWL<443> A_IWL<442> A_IWL<441> A_IWL<440> A_IWL<439> A_IWL<438> A_IWL<437> A_IWL<436> A_IWL<435> A_IWL<434> A_IWL<433> A_IWL<432> A_IWL<431> A_IWL<430> A_IWL<429> A_IWL<428> A_IWL<427> A_IWL<426> A_IWL<425> A_IWL<424> A_IWL<423> A_IWL<422> A_IWL<421> A_IWL<420> A_IWL<419> A_IWL<418> A_IWL<417> A_IWL<416> A_IWL<415> A_IWL<414> A_IWL<413> A_IWL<412> A_IWL<411> A_IWL<410> A_IWL<409> A_IWL<408> A_IWL<407> A_IWL<406> A_IWL<405> A_IWL<404> A_IWL<403> A_IWL<402> A_IWL<401> A_IWL<400> A_IWL<399> A_IWL<398> A_IWL<397> A_IWL<396> A_IWL<395> A_IWL<394> A_IWL<393> A_IWL<392> A_IWL<391> A_IWL<390> A_IWL<389> A_IWL<388> A_IWL<387> A_IWL<386> A_IWL<385> A_IWL<384> A_IWL<383> A_IWL<382> A_IWL<381> A_IWL<380> A_IWL<379> A_IWL<378> A_IWL<377> A_IWL<376> A_IWL<375> A_IWL<374> A_IWL<373> A_IWL<372> A_IWL<371> A_IWL<370> A_IWL<369> A_IWL<368> A_IWL<367> A_IWL<366> A_IWL<365> A_IWL<364> A_IWL<363> A_IWL<362> A_IWL<361> A_IWL<360> A_IWL<359> A_IWL<358> A_IWL<357> A_IWL<356> A_IWL<355> A_IWL<354> A_IWL<353> A_IWL<352> A_IWL<351> A_IWL<350> A_IWL<349> A_IWL<348> A_IWL<347> A_IWL<346> A_IWL<345> A_IWL<344> A_IWL<343> A_IWL<342> A_IWL<341> A_IWL<340> A_IWL<339> A_IWL<338> A_IWL<337> A_IWL<336> A_IWL<335> A_IWL<334> A_IWL<333> A_IWL<332> A_IWL<331> A_IWL<330> A_IWL<329> A_IWL<328> A_IWL<327> A_IWL<326> A_IWL<325> A_IWL<324> A_IWL<323> A_IWL<322> A_IWL<321> A_IWL<320> A_IWL<319> A_IWL<318> A_IWL<317> A_IWL<316> A_IWL<315> A_IWL<314> A_IWL<313> A_IWL<312> A_IWL<311> A_IWL<310> A_IWL<309> A_IWL<308> A_IWL<307> A_IWL<306> A_IWL<305> A_IWL<304> A_IWL<303> A_IWL<302> A_IWL<301> A_IWL<300> A_IWL<299> A_IWL<298> A_IWL<297> A_IWL<296> A_IWL<295> A_IWL<294> A_IWL<293> A_IWL<292> A_IWL<291> A_IWL<290> A_IWL<289> A_IWL<288> A_IWL<287> A_IWL<286> A_IWL<285> A_IWL<284> A_IWL<283> A_IWL<282> A_IWL<281> A_IWL<280> A_IWL<279> A_IWL<278> A_IWL<277> A_IWL<276> A_IWL<275> A_IWL<274> A_IWL<273> A_IWL<272> A_IWL<271> A_IWL<270> A_IWL<269> A_IWL<268> A_IWL<267> A_IWL<266> A_IWL<265> A_IWL<264> A_IWL<263> A_IWL<262> A_IWL<261> A_IWL<260> A_IWL<259> A_IWL<258> A_IWL<257> A_IWL<256> A_IWL<767> A_IWL<766> A_IWL<765> A_IWL<764> A_IWL<763> A_IWL<762> A_IWL<761> A_IWL<760> A_IWL<759> A_IWL<758> A_IWL<757> A_IWL<756> A_IWL<755> A_IWL<754> A_IWL<753> A_IWL<752> A_IWL<751> A_IWL<750> A_IWL<749> A_IWL<748> A_IWL<747> A_IWL<746> A_IWL<745> A_IWL<744> A_IWL<743> A_IWL<742> A_IWL<741> A_IWL<740> A_IWL<739> A_IWL<738> A_IWL<737> A_IWL<736> A_IWL<735> A_IWL<734> A_IWL<733> A_IWL<732> A_IWL<731> A_IWL<730> A_IWL<729> A_IWL<728> A_IWL<727> A_IWL<726> A_IWL<725> A_IWL<724> A_IWL<723> A_IWL<722> A_IWL<721> A_IWL<720> A_IWL<719> A_IWL<718> A_IWL<717> A_IWL<716> A_IWL<715> A_IWL<714> A_IWL<713> A_IWL<712> A_IWL<711> A_IWL<710> A_IWL<709> A_IWL<708> A_IWL<707> A_IWL<706> A_IWL<705> A_IWL<704> A_IWL<703> A_IWL<702> A_IWL<701> A_IWL<700> A_IWL<699> A_IWL<698> A_IWL<697> A_IWL<696> A_IWL<695> A_IWL<694> A_IWL<693> A_IWL<692> A_IWL<691> A_IWL<690> A_IWL<689> A_IWL<688> A_IWL<687> A_IWL<686> A_IWL<685> A_IWL<684> A_IWL<683> A_IWL<682> A_IWL<681> A_IWL<680> A_IWL<679> A_IWL<678> A_IWL<677> A_IWL<676> A_IWL<675> A_IWL<674> A_IWL<673> A_IWL<672> A_IWL<671> A_IWL<670> A_IWL<669> A_IWL<668> A_IWL<667> A_IWL<666> A_IWL<665> A_IWL<664> A_IWL<663> A_IWL<662> A_IWL<661> A_IWL<660> A_IWL<659> A_IWL<658> A_IWL<657> A_IWL<656> A_IWL<655> A_IWL<654> A_IWL<653> A_IWL<652> A_IWL<651> A_IWL<650> A_IWL<649> A_IWL<648> A_IWL<647> A_IWL<646> A_IWL<645> A_IWL<644> A_IWL<643> A_IWL<642> A_IWL<641> A_IWL<640> A_IWL<639> A_IWL<638> A_IWL<637> A_IWL<636> A_IWL<635> A_IWL<634> A_IWL<633> A_IWL<632> A_IWL<631> A_IWL<630> A_IWL<629> A_IWL<628> A_IWL<627> A_IWL<626> A_IWL<625> A_IWL<624> A_IWL<623> A_IWL<622> A_IWL<621> A_IWL<620> A_IWL<619> A_IWL<618> A_IWL<617> A_IWL<616> A_IWL<615> A_IWL<614> A_IWL<613> A_IWL<612> A_IWL<611> A_IWL<610> A_IWL<609> A_IWL<608> A_IWL<607> A_IWL<606> A_IWL<605> A_IWL<604> A_IWL<603> A_IWL<602> A_IWL<601> A_IWL<600> A_IWL<599> A_IWL<598> A_IWL<597> A_IWL<596> A_IWL<595> A_IWL<594> A_IWL<593> A_IWL<592> A_IWL<591> A_IWL<590> A_IWL<589> A_IWL<588> A_IWL<587> A_IWL<586> A_IWL<585> A_IWL<584> A_IWL<583> A_IWL<582> A_IWL<581> A_IWL<580> A_IWL<579> A_IWL<578> A_IWL<577> A_IWL<576> A_IWL<575> A_IWL<574> A_IWL<573> A_IWL<572> A_IWL<571> A_IWL<570> A_IWL<569> A_IWL<568> A_IWL<567> A_IWL<566> A_IWL<565> A_IWL<564> A_IWL<563> A_IWL<562> A_IWL<561> A_IWL<560> A_IWL<559> A_IWL<558> A_IWL<557> A_IWL<556> A_IWL<555> A_IWL<554> A_IWL<553> A_IWL<552> A_IWL<551> A_IWL<550> A_IWL<549> A_IWL<548> A_IWL<547> A_IWL<546> A_IWL<545> A_IWL<544> A_IWL<543> A_IWL<542> A_IWL<541> A_IWL<540> A_IWL<539> A_IWL<538> A_IWL<537> A_IWL<536> A_IWL<535> A_IWL<534> A_IWL<533> A_IWL<532> A_IWL<531> A_IWL<530> A_IWL<529> A_IWL<528> A_IWL<527> A_IWL<526> A_IWL<525> A_IWL<524> A_IWL<523> A_IWL<522> A_IWL<521> A_IWL<520> A_IWL<519> A_IWL<518> A_IWL<517> A_IWL<516> A_IWL<515> A_IWL<514> A_IWL<513> A_IWL<512> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<1> A_BLC<3> A_BLC<2> A_BLC_TOP<3> A_BLC_TOP<2> A_BLT<3> A_BLT<2> A_BLT_TOP<3> A_BLT_TOP<2> A_IWL<255> A_IWL<254> A_IWL<253> A_IWL<252> A_IWL<251> A_IWL<250> A_IWL<249> A_IWL<248> A_IWL<247> A_IWL<246> A_IWL<245> A_IWL<244> A_IWL<243> A_IWL<242> A_IWL<241> A_IWL<240> A_IWL<239> A_IWL<238> A_IWL<237> A_IWL<236> A_IWL<235> A_IWL<234> A_IWL<233> A_IWL<232> A_IWL<231> A_IWL<230> A_IWL<229> A_IWL<228> A_IWL<227> A_IWL<226> A_IWL<225> A_IWL<224> A_IWL<223> A_IWL<222> A_IWL<221> A_IWL<220> A_IWL<219> A_IWL<218> A_IWL<217> A_IWL<216> A_IWL<215> A_IWL<214> A_IWL<213> A_IWL<212> A_IWL<211> A_IWL<210> A_IWL<209> A_IWL<208> A_IWL<207> A_IWL<206> A_IWL<205> A_IWL<204> A_IWL<203> A_IWL<202> A_IWL<201> A_IWL<200> A_IWL<199> A_IWL<198> A_IWL<197> A_IWL<196> A_IWL<195> A_IWL<194> A_IWL<193> A_IWL<192> A_IWL<191> A_IWL<190> A_IWL<189> A_IWL<188> A_IWL<187> A_IWL<186> A_IWL<185> A_IWL<184> A_IWL<183> A_IWL<182> A_IWL<181> A_IWL<180> A_IWL<179> A_IWL<178> A_IWL<177> A_IWL<176> A_IWL<175> A_IWL<174> A_IWL<173> A_IWL<172> A_IWL<171> A_IWL<170> A_IWL<169> A_IWL<168> A_IWL<167> A_IWL<166> A_IWL<165> A_IWL<164> A_IWL<163> A_IWL<162> A_IWL<161> A_IWL<160> A_IWL<159> A_IWL<158> A_IWL<157> A_IWL<156> A_IWL<155> A_IWL<154> A_IWL<153> A_IWL<152> A_IWL<151> A_IWL<150> A_IWL<149> A_IWL<148> A_IWL<147> A_IWL<146> A_IWL<145> A_IWL<144> A_IWL<143> A_IWL<142> A_IWL<141> A_IWL<140> A_IWL<139> A_IWL<138> A_IWL<137> A_IWL<136> A_IWL<135> A_IWL<134> A_IWL<133> A_IWL<132> A_IWL<131> A_IWL<130> A_IWL<129> A_IWL<128> A_IWL<127> A_IWL<126> A_IWL<125> A_IWL<124> A_IWL<123> A_IWL<122> A_IWL<121> A_IWL<120> A_IWL<119> A_IWL<118> A_IWL<117> A_IWL<116> A_IWL<115> A_IWL<114> A_IWL<113> A_IWL<112> A_IWL<111> A_IWL<110> A_IWL<109> A_IWL<108> A_IWL<107> A_IWL<106> A_IWL<105> A_IWL<104> A_IWL<103> A_IWL<102> A_IWL<101> A_IWL<100> A_IWL<99> A_IWL<98> A_IWL<97> A_IWL<96> A_IWL<95> A_IWL<94> A_IWL<93> A_IWL<92> A_IWL<91> A_IWL<90> A_IWL<89> A_IWL<88> A_IWL<87> A_IWL<86> A_IWL<85> A_IWL<84> A_IWL<83> A_IWL<82> A_IWL<81> A_IWL<80> A_IWL<79> A_IWL<78> A_IWL<77> A_IWL<76> A_IWL<75> A_IWL<74> A_IWL<73> A_IWL<72> A_IWL<71> A_IWL<70> A_IWL<69> A_IWL<68> A_IWL<67> A_IWL<66> A_IWL<65> A_IWL<64> A_IWL<63> A_IWL<62> A_IWL<61> A_IWL<60> A_IWL<59> A_IWL<58> A_IWL<57> A_IWL<56> A_IWL<55> A_IWL<54> A_IWL<53> A_IWL<52> A_IWL<51> A_IWL<50> A_IWL<49> A_IWL<48> A_IWL<47> A_IWL<46> A_IWL<45> A_IWL<44> A_IWL<43> A_IWL<42> A_IWL<41> A_IWL<40> A_IWL<39> A_IWL<38> A_IWL<37> A_IWL<36> A_IWL<35> A_IWL<34> A_IWL<33> A_IWL<32> A_IWL<31> A_IWL<30> A_IWL<29> A_IWL<28> A_IWL<27> A_IWL<26> A_IWL<25> A_IWL<24> A_IWL<23> A_IWL<22> A_IWL<21> A_IWL<20> A_IWL<19> A_IWL<18> A_IWL<17> A_IWL<16> A_IWL<15> A_IWL<14> A_IWL<13> A_IWL<12> A_IWL<11> A_IWL<10> A_IWL<9> A_IWL<8> A_IWL<7> A_IWL<6> A_IWL<5> A_IWL<4> A_IWL<3> A_IWL<2> A_IWL<1> A_IWL<0> A_IWL<511> A_IWL<510> A_IWL<509> A_IWL<508> A_IWL<507> A_IWL<506> A_IWL<505> A_IWL<504> A_IWL<503> A_IWL<502> A_IWL<501> A_IWL<500> A_IWL<499> A_IWL<498> A_IWL<497> A_IWL<496> A_IWL<495> A_IWL<494> A_IWL<493> A_IWL<492> A_IWL<491> A_IWL<490> A_IWL<489> A_IWL<488> A_IWL<487> A_IWL<486> A_IWL<485> A_IWL<484> A_IWL<483> A_IWL<482> A_IWL<481> A_IWL<480> A_IWL<479> A_IWL<478> A_IWL<477> A_IWL<476> A_IWL<475> A_IWL<474> A_IWL<473> A_IWL<472> A_IWL<471> A_IWL<470> A_IWL<469> A_IWL<468> A_IWL<467> A_IWL<466> A_IWL<465> A_IWL<464> A_IWL<463> A_IWL<462> A_IWL<461> A_IWL<460> A_IWL<459> A_IWL<458> A_IWL<457> A_IWL<456> A_IWL<455> A_IWL<454> A_IWL<453> A_IWL<452> A_IWL<451> A_IWL<450> A_IWL<449> A_IWL<448> A_IWL<447> A_IWL<446> A_IWL<445> A_IWL<444> A_IWL<443> A_IWL<442> A_IWL<441> A_IWL<440> A_IWL<439> A_IWL<438> A_IWL<437> A_IWL<436> A_IWL<435> A_IWL<434> A_IWL<433> A_IWL<432> A_IWL<431> A_IWL<430> A_IWL<429> A_IWL<428> A_IWL<427> A_IWL<426> A_IWL<425> A_IWL<424> A_IWL<423> A_IWL<422> A_IWL<421> A_IWL<420> A_IWL<419> A_IWL<418> A_IWL<417> A_IWL<416> A_IWL<415> A_IWL<414> A_IWL<413> A_IWL<412> A_IWL<411> A_IWL<410> A_IWL<409> A_IWL<408> A_IWL<407> A_IWL<406> A_IWL<405> A_IWL<404> A_IWL<403> A_IWL<402> A_IWL<401> A_IWL<400> A_IWL<399> A_IWL<398> A_IWL<397> A_IWL<396> A_IWL<395> A_IWL<394> A_IWL<393> A_IWL<392> A_IWL<391> A_IWL<390> A_IWL<389> A_IWL<388> A_IWL<387> A_IWL<386> A_IWL<385> A_IWL<384> A_IWL<383> A_IWL<382> A_IWL<381> A_IWL<380> A_IWL<379> A_IWL<378> A_IWL<377> A_IWL<376> A_IWL<375> A_IWL<374> A_IWL<373> A_IWL<372> A_IWL<371> A_IWL<370> A_IWL<369> A_IWL<368> A_IWL<367> A_IWL<366> A_IWL<365> A_IWL<364> A_IWL<363> A_IWL<362> A_IWL<361> A_IWL<360> A_IWL<359> A_IWL<358> A_IWL<357> A_IWL<356> A_IWL<355> A_IWL<354> A_IWL<353> A_IWL<352> A_IWL<351> A_IWL<350> A_IWL<349> A_IWL<348> A_IWL<347> A_IWL<346> A_IWL<345> A_IWL<344> A_IWL<343> A_IWL<342> A_IWL<341> A_IWL<340> A_IWL<339> A_IWL<338> A_IWL<337> A_IWL<336> A_IWL<335> A_IWL<334> A_IWL<333> A_IWL<332> A_IWL<331> A_IWL<330> A_IWL<329> A_IWL<328> A_IWL<327> A_IWL<326> A_IWL<325> A_IWL<324> A_IWL<323> A_IWL<322> A_IWL<321> A_IWL<320> A_IWL<319> A_IWL<318> A_IWL<317> A_IWL<316> A_IWL<315> A_IWL<314> A_IWL<313> A_IWL<312> A_IWL<311> A_IWL<310> A_IWL<309> A_IWL<308> A_IWL<307> A_IWL<306> A_IWL<305> A_IWL<304> A_IWL<303> A_IWL<302> A_IWL<301> A_IWL<300> A_IWL<299> A_IWL<298> A_IWL<297> A_IWL<296> A_IWL<295> A_IWL<294> A_IWL<293> A_IWL<292> A_IWL<291> A_IWL<290> A_IWL<289> A_IWL<288> A_IWL<287> A_IWL<286> A_IWL<285> A_IWL<284> A_IWL<283> A_IWL<282> A_IWL<281> A_IWL<280> A_IWL<279> A_IWL<278> A_IWL<277> A_IWL<276> A_IWL<275> A_IWL<274> A_IWL<273> A_IWL<272> A_IWL<271> A_IWL<270> A_IWL<269> A_IWL<268> A_IWL<267> A_IWL<266> A_IWL<265> A_IWL<264> A_IWL<263> A_IWL<262> A_IWL<261> A_IWL<260> A_IWL<259> A_IWL<258> A_IWL<257> A_IWL<256> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
XCOL<0> A_BLC<1> A_BLC<0> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT<1> A_BLT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_WL<255> A_WL<254> A_WL<253> A_WL<252> A_WL<251> A_WL<250> A_WL<249> A_WL<248> A_WL<247> A_WL<246> A_WL<245> A_WL<244> A_WL<243> A_WL<242> A_WL<241> A_WL<240> A_WL<239> A_WL<238> A_WL<237> A_WL<236> A_WL<235> A_WL<234> A_WL<233> A_WL<232> A_WL<231> A_WL<230> A_WL<229> A_WL<228> A_WL<227> A_WL<226> A_WL<225> A_WL<224> A_WL<223> A_WL<222> A_WL<221> A_WL<220> A_WL<219> A_WL<218> A_WL<217> A_WL<216> A_WL<215> A_WL<214> A_WL<213> A_WL<212> A_WL<211> A_WL<210> A_WL<209> A_WL<208> A_WL<207> A_WL<206> A_WL<205> A_WL<204> A_WL<203> A_WL<202> A_WL<201> A_WL<200> A_WL<199> A_WL<198> A_WL<197> A_WL<196> A_WL<195> A_WL<194> A_WL<193> A_WL<192> A_WL<191> A_WL<190> A_WL<189> A_WL<188> A_WL<187> A_WL<186> A_WL<185> A_WL<184> A_WL<183> A_WL<182> A_WL<181> A_WL<180> A_WL<179> A_WL<178> A_WL<177> A_WL<176> A_WL<175> A_WL<174> A_WL<173> A_WL<172> A_WL<171> A_WL<170> A_WL<169> A_WL<168> A_WL<167> A_WL<166> A_WL<165> A_WL<164> A_WL<163> A_WL<162> A_WL<161> A_WL<160> A_WL<159> A_WL<158> A_WL<157> A_WL<156> A_WL<155> A_WL<154> A_WL<153> A_WL<152> A_WL<151> A_WL<150> A_WL<149> A_WL<148> A_WL<147> A_WL<146> A_WL<145> A_WL<144> A_WL<143> A_WL<142> A_WL<141> A_WL<140> A_WL<139> A_WL<138> A_WL<137> A_WL<136> A_WL<135> A_WL<134> A_WL<133> A_WL<132> A_WL<131> A_WL<130> A_WL<129> A_WL<128> A_WL<127> A_WL<126> A_WL<125> A_WL<124> A_WL<123> A_WL<122> A_WL<121> A_WL<120> A_WL<119> A_WL<118> A_WL<117> A_WL<116> A_WL<115> A_WL<114> A_WL<113> A_WL<112> A_WL<111> A_WL<110> A_WL<109> A_WL<108> A_WL<107> A_WL<106> A_WL<105> A_WL<104> A_WL<103> A_WL<102> A_WL<101> A_WL<100> A_WL<99> A_WL<98> A_WL<97> A_WL<96> A_WL<95> A_WL<94> A_WL<93> A_WL<92> A_WL<91> A_WL<90> A_WL<89> A_WL<88> A_WL<87> A_WL<86> A_WL<85> A_WL<84> A_WL<83> A_WL<82> A_WL<81> A_WL<80> A_WL<79> A_WL<78> A_WL<77> A_WL<76> A_WL<75> A_WL<74> A_WL<73> A_WL<72> A_WL<71> A_WL<70> A_WL<69> A_WL<68> A_WL<67> A_WL<66> A_WL<65> A_WL<64> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> A_IWL<255> A_IWL<254> A_IWL<253> A_IWL<252> A_IWL<251> A_IWL<250> A_IWL<249> A_IWL<248> A_IWL<247> A_IWL<246> A_IWL<245> A_IWL<244> A_IWL<243> A_IWL<242> A_IWL<241> A_IWL<240> A_IWL<239> A_IWL<238> A_IWL<237> A_IWL<236> A_IWL<235> A_IWL<234> A_IWL<233> A_IWL<232> A_IWL<231> A_IWL<230> A_IWL<229> A_IWL<228> A_IWL<227> A_IWL<226> A_IWL<225> A_IWL<224> A_IWL<223> A_IWL<222> A_IWL<221> A_IWL<220> A_IWL<219> A_IWL<218> A_IWL<217> A_IWL<216> A_IWL<215> A_IWL<214> A_IWL<213> A_IWL<212> A_IWL<211> A_IWL<210> A_IWL<209> A_IWL<208> A_IWL<207> A_IWL<206> A_IWL<205> A_IWL<204> A_IWL<203> A_IWL<202> A_IWL<201> A_IWL<200> A_IWL<199> A_IWL<198> A_IWL<197> A_IWL<196> A_IWL<195> A_IWL<194> A_IWL<193> A_IWL<192> A_IWL<191> A_IWL<190> A_IWL<189> A_IWL<188> A_IWL<187> A_IWL<186> A_IWL<185> A_IWL<184> A_IWL<183> A_IWL<182> A_IWL<181> A_IWL<180> A_IWL<179> A_IWL<178> A_IWL<177> A_IWL<176> A_IWL<175> A_IWL<174> A_IWL<173> A_IWL<172> A_IWL<171> A_IWL<170> A_IWL<169> A_IWL<168> A_IWL<167> A_IWL<166> A_IWL<165> A_IWL<164> A_IWL<163> A_IWL<162> A_IWL<161> A_IWL<160> A_IWL<159> A_IWL<158> A_IWL<157> A_IWL<156> A_IWL<155> A_IWL<154> A_IWL<153> A_IWL<152> A_IWL<151> A_IWL<150> A_IWL<149> A_IWL<148> A_IWL<147> A_IWL<146> A_IWL<145> A_IWL<144> A_IWL<143> A_IWL<142> A_IWL<141> A_IWL<140> A_IWL<139> A_IWL<138> A_IWL<137> A_IWL<136> A_IWL<135> A_IWL<134> A_IWL<133> A_IWL<132> A_IWL<131> A_IWL<130> A_IWL<129> A_IWL<128> A_IWL<127> A_IWL<126> A_IWL<125> A_IWL<124> A_IWL<123> A_IWL<122> A_IWL<121> A_IWL<120> A_IWL<119> A_IWL<118> A_IWL<117> A_IWL<116> A_IWL<115> A_IWL<114> A_IWL<113> A_IWL<112> A_IWL<111> A_IWL<110> A_IWL<109> A_IWL<108> A_IWL<107> A_IWL<106> A_IWL<105> A_IWL<104> A_IWL<103> A_IWL<102> A_IWL<101> A_IWL<100> A_IWL<99> A_IWL<98> A_IWL<97> A_IWL<96> A_IWL<95> A_IWL<94> A_IWL<93> A_IWL<92> A_IWL<91> A_IWL<90> A_IWL<89> A_IWL<88> A_IWL<87> A_IWL<86> A_IWL<85> A_IWL<84> A_IWL<83> A_IWL<82> A_IWL<81> A_IWL<80> A_IWL<79> A_IWL<78> A_IWL<77> A_IWL<76> A_IWL<75> A_IWL<74> A_IWL<73> A_IWL<72> A_IWL<71> A_IWL<70> A_IWL<69> A_IWL<68> A_IWL<67> A_IWL<66> A_IWL<65> A_IWL<64> A_IWL<63> A_IWL<62> A_IWL<61> A_IWL<60> A_IWL<59> A_IWL<58> A_IWL<57> A_IWL<56> A_IWL<55> A_IWL<54> A_IWL<53> A_IWL<52> A_IWL<51> A_IWL<50> A_IWL<49> A_IWL<48> A_IWL<47> A_IWL<46> A_IWL<45> A_IWL<44> A_IWL<43> A_IWL<42> A_IWL<41> A_IWL<40> A_IWL<39> A_IWL<38> A_IWL<37> A_IWL<36> A_IWL<35> A_IWL<34> A_IWL<33> A_IWL<32> A_IWL<31> A_IWL<30> A_IWL<29> A_IWL<28> A_IWL<27> A_IWL<26> A_IWL<25> A_IWL<24> A_IWL<23> A_IWL<22> A_IWL<21> A_IWL<20> A_IWL<19> A_IWL<18> A_IWL<17> A_IWL<16> A_IWL<15> A_IWL<14> A_IWL<13> A_IWL<12> A_IWL<11> A_IWL<10> A_IWL<9> A_IWL<8> A_IWL<7> A_IWL<6> A_IWL<5> A_IWL<4> A_IWL<3> A_IWL<2> A_IWL<1> A_IWL<0> VDD_CORE VSS / RM_IHPSG13_1024x64_c2_1P_COLUMN_pcell_0
.ENDS




.SUBCKT RM_IHPSG13_1024x64_c2_1P_DLY_pcell_2 A Z VDD VSS
	XIDL<2> D<7> Z VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<1> D<6> D<7> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDM<6> D<5> D<6> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<5> D<4> D<5> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<4> D<3> D<4> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
.ENDS


.SUBCKT RM_IHPSG13_1024x64_c2_1P_DLY_pcell_3 A Z VDD VSS
	XIDL<4> D<7> Z VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<3> D<6> D<7> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<2> D<5> D<6> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<1> D<4> D<5> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDM<4> D<3> D<4> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
.ENDS



.SUBCKT RM_IHPSG13_1P_1024x64_c2_bm_bist A_ADDR<9> A_ADDR<8> A_ADDR<7> A_ADDR<6> A_ADDR<5> A_ADDR<4> A_ADDR<3> A_ADDR<2> A_ADDR<1> A_ADDR<0> A_BIST_ADDR<9> A_BIST_ADDR<8> A_BIST_ADDR<7> A_BIST_ADDR<6> A_BIST_ADDR<5> A_BIST_ADDR<4> A_BIST_ADDR<3> A_BIST_ADDR<2> A_BIST_ADDR<1> A_BIST_ADDR<0> A_BIST_BM<63> A_BIST_BM<62> A_BIST_BM<61> A_BIST_BM<60> A_BIST_BM<59> A_BIST_BM<58> A_BIST_BM<57> A_BIST_BM<56> A_BIST_BM<55> A_BIST_BM<54> A_BIST_BM<53> A_BIST_BM<52> A_BIST_BM<51> A_BIST_BM<50> A_BIST_BM<49> A_BIST_BM<48> A_BIST_BM<47> A_BIST_BM<46> A_BIST_BM<45> A_BIST_BM<44> A_BIST_BM<43> A_BIST_BM<42> A_BIST_BM<41> A_BIST_BM<40> A_BIST_BM<39> A_BIST_BM<38> A_BIST_BM<37> A_BIST_BM<36> A_BIST_BM<35> A_BIST_BM<34> A_BIST_BM<33> A_BIST_BM<32> A_BIST_BM<31> A_BIST_BM<30> A_BIST_BM<29> A_BIST_BM<28> A_BIST_BM<27> A_BIST_BM<26> A_BIST_BM<25> A_BIST_BM<24> A_BIST_BM<23> A_BIST_BM<22> A_BIST_BM<21> A_BIST_BM<20> A_BIST_BM<19> A_BIST_BM<18> A_BIST_BM<17> A_BIST_BM<16> A_BIST_BM<15> A_BIST_BM<14> A_BIST_BM<13> A_BIST_BM<12> A_BIST_BM<11> A_BIST_BM<10> A_BIST_BM<9> A_BIST_BM<8> A_BIST_BM<7> A_BIST_BM<6> A_BIST_BM<5> A_BIST_BM<4> A_BIST_BM<3> A_BIST_BM<2> A_BIST_BM<1> A_BIST_BM<0> A_BIST_CLK A_BIST_DIN<63> A_BIST_DIN<62> A_BIST_DIN<61> A_BIST_DIN<60> A_BIST_DIN<59> A_BIST_DIN<58> A_BIST_DIN<57> A_BIST_DIN<56> A_BIST_DIN<55> A_BIST_DIN<54> A_BIST_DIN<53> A_BIST_DIN<52> A_BIST_DIN<51> A_BIST_DIN<50> A_BIST_DIN<49> A_BIST_DIN<48> A_BIST_DIN<47> A_BIST_DIN<46> A_BIST_DIN<45> A_BIST_DIN<44> A_BIST_DIN<43> A_BIST_DIN<42> A_BIST_DIN<41> A_BIST_DIN<40> A_BIST_DIN<39> A_BIST_DIN<38> A_BIST_DIN<37> A_BIST_DIN<36> A_BIST_DIN<35> A_BIST_DIN<34> A_BIST_DIN<33> A_BIST_DIN<32> A_BIST_DIN<31> A_BIST_DIN<30> A_BIST_DIN<29> A_BIST_DIN<28> A_BIST_DIN<27> A_BIST_DIN<26> A_BIST_DIN<25> A_BIST_DIN<24> A_BIST_DIN<23> A_BIST_DIN<22> A_BIST_DIN<21> A_BIST_DIN<20> A_BIST_DIN<19> A_BIST_DIN<18> A_BIST_DIN<17> A_BIST_DIN<16> A_BIST_DIN<15> A_BIST_DIN<14> A_BIST_DIN<13> A_BIST_DIN<12> A_BIST_DIN<11> A_BIST_DIN<10> A_BIST_DIN<9> A_BIST_DIN<8> A_BIST_DIN<7> A_BIST_DIN<6> A_BIST_DIN<5> A_BIST_DIN<4> A_BIST_DIN<3> A_BIST_DIN<2> A_BIST_DIN<1> A_BIST_DIN<0> A_BIST_EN A_BIST_MEN A_BIST_REN A_BIST_WEN A_BM<63> A_BM<62> A_BM<61> A_BM<60> A_BM<59> A_BM<58> A_BM<57> A_BM<56> A_BM<55> A_BM<54> A_BM<53> A_BM<52> A_BM<51> A_BM<50> A_BM<49> A_BM<48> A_BM<47> A_BM<46> A_BM<45> A_BM<44> A_BM<43> A_BM<42> A_BM<41> A_BM<40> A_BM<39> A_BM<38> A_BM<37> A_BM<36> A_BM<35> A_BM<34> A_BM<33> A_BM<32> A_BM<31> A_BM<30> A_BM<29> A_BM<28> A_BM<27> A_BM<26> A_BM<25> A_BM<24> A_BM<23> A_BM<22> A_BM<21> A_BM<20> A_BM<19> A_BM<18> A_BM<17> A_BM<16> A_BM<15> A_BM<14> A_BM<13> A_BM<12> A_BM<11> A_BM<10> A_BM<9> A_BM<8> A_BM<7> A_BM<6> A_BM<5> A_BM<4> A_BM<3> A_BM<2> A_BM<1> A_BM<0> A_CLK A_DIN<63> A_DIN<62> A_DIN<61> A_DIN<60> A_DIN<59> A_DIN<58> A_DIN<57> A_DIN<56> A_DIN<55> A_DIN<54> A_DIN<53> A_DIN<52> A_DIN<51> A_DIN<50> A_DIN<49> A_DIN<48> A_DIN<47> A_DIN<46> A_DIN<45> A_DIN<44> A_DIN<43> A_DIN<42> A_DIN<41> A_DIN<40> A_DIN<39> A_DIN<38> A_DIN<37> A_DIN<36> A_DIN<35> A_DIN<34> A_DIN<33> A_DIN<32> A_DIN<31> A_DIN<30> A_DIN<29> A_DIN<28> A_DIN<27> A_DIN<26> A_DIN<25> A_DIN<24> A_DIN<23> A_DIN<22> A_DIN<21> A_DIN<20> A_DIN<19> A_DIN<18> A_DIN<17> A_DIN<16> A_DIN<15> A_DIN<14> A_DIN<13> A_DIN<12> A_DIN<11> A_DIN<10> A_DIN<9> A_DIN<8> A_DIN<7> A_DIN<6> A_DIN<5> A_DIN<4> A_DIN<3> A_DIN<2> A_DIN<1> A_DIN<0> A_DLY A_DOUT<63> A_DOUT<62> A_DOUT<61> A_DOUT<60> A_DOUT<59> A_DOUT<58> A_DOUT<57> A_DOUT<56> A_DOUT<55> A_DOUT<54> A_DOUT<53> A_DOUT<52> A_DOUT<51> A_DOUT<50> A_DOUT<49> A_DOUT<48> A_DOUT<47> A_DOUT<46> A_DOUT<45> A_DOUT<44> A_DOUT<43> A_DOUT<42> A_DOUT<41> A_DOUT<40> A_DOUT<39> A_DOUT<38> A_DOUT<37> A_DOUT<36> A_DOUT<35> A_DOUT<34> A_DOUT<33> A_DOUT<32> A_DOUT<31> A_DOUT<30> A_DOUT<29> A_DOUT<28> A_DOUT<27> A_DOUT<26> A_DOUT<25> A_DOUT<24> A_DOUT<23> A_DOUT<22> A_DOUT<21> A_DOUT<20> A_DOUT<19> A_DOUT<18> A_DOUT<17> A_DOUT<16> A_DOUT<15> A_DOUT<14> A_DOUT<13> A_DOUT<12> A_DOUT<11> A_DOUT<10> A_DOUT<9> A_DOUT<8> A_DOUT<7> A_DOUT<6> A_DOUT<5> A_DOUT<4> A_DOUT<3> A_DOUT<2> A_DOUT<1> A_DOUT<0> A_MEN A_REN A_WEN VDD! VDDARRAY! VSS!


XRAM<1> a_blc_r<127> a_blc_r<126> a_blc_r<125> a_blc_r<124> a_blc_r<123> a_blc_r<122> a_blc_r<121> a_blc_r<120> a_blc_r<119> a_blc_r<118> a_blc_r<117> a_blc_r<116> a_blc_r<115> a_blc_r<114> a_blc_r<113> a_blc_r<112> a_blc_r<111> a_blc_r<110> a_blc_r<109> a_blc_r<108> a_blc_r<107> a_blc_r<106> a_blc_r<105> a_blc_r<104> a_blc_r<103> a_blc_r<102> a_blc_r<101> a_blc_r<100> a_blc_r<99> a_blc_r<98> a_blc_r<97> a_blc_r<96> a_blc_r<95> a_blc_r<94> a_blc_r<93> a_blc_r<92> a_blc_r<91> a_blc_r<90> a_blc_r<89> a_blc_r<88> a_blc_r<87> a_blc_r<86> a_blc_r<85> a_blc_r<84> a_blc_r<83> a_blc_r<82> a_blc_r<81> a_blc_r<80> a_blc_r<79> a_blc_r<78> a_blc_r<77> a_blc_r<76> a_blc_r<75> a_blc_r<74> a_blc_r<73> a_blc_r<72> a_blc_r<71> a_blc_r<70> a_blc_r<69> a_blc_r<68> a_blc_r<67> a_blc_r<66> a_blc_r<65> a_blc_r<64> a_blc_r<63> a_blc_r<62> a_blc_r<61> a_blc_r<60> a_blc_r<59> a_blc_r<58> a_blc_r<57> a_blc_r<56> a_blc_r<55> a_blc_r<54> a_blc_r<53> a_blc_r<52> a_blc_r<51> a_blc_r<50> a_blc_r<49> a_blc_r<48> a_blc_r<47> a_blc_r<46> a_blc_r<45> a_blc_r<44> a_blc_r<43> a_blc_r<42> a_blc_r<41> a_blc_r<40> a_blc_r<39> a_blc_r<38> a_blc_r<37> a_blc_r<36> a_blc_r<35> a_blc_r<34> a_blc_r<33> a_blc_r<32> a_blc_r<31> a_blc_r<30> a_blc_r<29> a_blc_r<28> a_blc_r<27> a_blc_r<26> a_blc_r<25> a_blc_r<24> a_blc_r<23> a_blc_r<22> a_blc_r<21> a_blc_r<20> a_blc_r<19> a_blc_r<18> a_blc_r<17> a_blc_r<16> a_blc_r<15> a_blc_r<14> a_blc_r<13> a_blc_r<12> a_blc_r<11> a_blc_r<10> a_blc_r<9> a_blc_r<8> a_blc_r<7> a_blc_r<6> a_blc_r<5> a_blc_r<4> a_blc_r<3> a_blc_r<2> a_blc_r<1> a_blc_r<0> a_blt_r<127> a_blt_r<126> a_blt_r<125> a_blt_r<124> a_blt_r<123> a_blt_r<122> a_blt_r<121> a_blt_r<120> a_blt_r<119> a_blt_r<118> a_blt_r<117> a_blt_r<116> a_blt_r<115> a_blt_r<114> a_blt_r<113> a_blt_r<112> a_blt_r<111> a_blt_r<110> a_blt_r<109> a_blt_r<108> a_blt_r<107> a_blt_r<106> a_blt_r<105> a_blt_r<104> a_blt_r<103> a_blt_r<102> a_blt_r<101> a_blt_r<100> a_blt_r<99> a_blt_r<98> a_blt_r<97> a_blt_r<96> a_blt_r<95> a_blt_r<94> a_blt_r<93> a_blt_r<92> a_blt_r<91> a_blt_r<90> a_blt_r<89> a_blt_r<88> a_blt_r<87> a_blt_r<86> a_blt_r<85> a_blt_r<84> a_blt_r<83> a_blt_r<82> a_blt_r<81> a_blt_r<80> a_blt_r<79> a_blt_r<78> a_blt_r<77> a_blt_r<76> a_blt_r<75> a_blt_r<74> a_blt_r<73> a_blt_r<72> a_blt_r<71> a_blt_r<70> a_blt_r<69> a_blt_r<68> a_blt_r<67> a_blt_r<66> a_blt_r<65> a_blt_r<64> a_blt_r<63> a_blt_r<62> a_blt_r<61> a_blt_r<60> a_blt_r<59> a_blt_r<58> a_blt_r<57> a_blt_r<56> a_blt_r<55> a_blt_r<54> a_blt_r<53> a_blt_r<52> a_blt_r<51> a_blt_r<50> a_blt_r<49> a_blt_r<48> a_blt_r<47> a_blt_r<46> a_blt_r<45> a_blt_r<44> a_blt_r<43> a_blt_r<42> a_blt_r<41> a_blt_r<40> a_blt_r<39> a_blt_r<38> a_blt_r<37> a_blt_r<36> a_blt_r<35> a_blt_r<34> a_blt_r<33> a_blt_r<32> a_blt_r<31> a_blt_r<30> a_blt_r<29> a_blt_r<28> a_blt_r<27> a_blt_r<26> a_blt_r<25> a_blt_r<24> a_blt_r<23> a_blt_r<22> a_blt_r<21> a_blt_r<20> a_blt_r<19> a_blt_r<18> a_blt_r<17> a_blt_r<16> a_blt_r<15> a_blt_r<14> a_blt_r<13> a_blt_r<12> a_blt_r<11> a_blt_r<10> a_blt_r<9> a_blt_r<8> a_blt_r<7> a_blt_r<6> a_blt_r<5> a_blt_r<4> a_blt_r<3> a_blt_r<2> a_blt_r<1> a_blt_r<0> a_wl_r<255> a_wl_r<254> a_wl_r<253> a_wl_r<252> a_wl_r<251> a_wl_r<250> a_wl_r<249> a_wl_r<248> a_wl_r<247> a_wl_r<246> a_wl_r<245> a_wl_r<244> a_wl_r<243> a_wl_r<242> a_wl_r<241> a_wl_r<240> a_wl_r<239> a_wl_r<238> a_wl_r<237> a_wl_r<236> a_wl_r<235> a_wl_r<234> a_wl_r<233> a_wl_r<232> a_wl_r<231> a_wl_r<230> a_wl_r<229> a_wl_r<228> a_wl_r<227> a_wl_r<226> a_wl_r<225> a_wl_r<224> a_wl_r<223> a_wl_r<222> a_wl_r<221> a_wl_r<220> a_wl_r<219> a_wl_r<218> a_wl_r<217> a_wl_r<216> a_wl_r<215> a_wl_r<214> a_wl_r<213> a_wl_r<212> a_wl_r<211> a_wl_r<210> a_wl_r<209> a_wl_r<208> a_wl_r<207> a_wl_r<206> a_wl_r<205> a_wl_r<204> a_wl_r<203> a_wl_r<202> a_wl_r<201> a_wl_r<200> a_wl_r<199> a_wl_r<198> a_wl_r<197> a_wl_r<196> a_wl_r<195> a_wl_r<194> a_wl_r<193> a_wl_r<192> a_wl_r<191> a_wl_r<190> a_wl_r<189> a_wl_r<188> a_wl_r<187> a_wl_r<186> a_wl_r<185> a_wl_r<184> a_wl_r<183> a_wl_r<182> a_wl_r<181> a_wl_r<180> a_wl_r<179> a_wl_r<178> a_wl_r<177> a_wl_r<176> a_wl_r<175> a_wl_r<174> a_wl_r<173> a_wl_r<172> a_wl_r<171> a_wl_r<170> a_wl_r<169> a_wl_r<168> a_wl_r<167> a_wl_r<166> a_wl_r<165> a_wl_r<164> a_wl_r<163> a_wl_r<162> a_wl_r<161> a_wl_r<160> a_wl_r<159> a_wl_r<158> a_wl_r<157> a_wl_r<156> a_wl_r<155> a_wl_r<154> a_wl_r<153> a_wl_r<152> a_wl_r<151> a_wl_r<150> a_wl_r<149> a_wl_r<148> a_wl_r<147> a_wl_r<146> a_wl_r<145> a_wl_r<144> a_wl_r<143> a_wl_r<142> a_wl_r<141> a_wl_r<140> a_wl_r<139> a_wl_r<138> a_wl_r<137> a_wl_r<136> a_wl_r<135> a_wl_r<134> a_wl_r<133> a_wl_r<132> a_wl_r<131> a_wl_r<130> a_wl_r<129> a_wl_r<128> a_wl_r<127> a_wl_r<126> a_wl_r<125> a_wl_r<124> a_wl_r<123> a_wl_r<122> a_wl_r<121> a_wl_r<120> a_wl_r<119> a_wl_r<118> a_wl_r<117> a_wl_r<116> a_wl_r<115> a_wl_r<114> a_wl_r<113> a_wl_r<112> a_wl_r<111> a_wl_r<110> a_wl_r<109> a_wl_r<108> a_wl_r<107> a_wl_r<106> a_wl_r<105> a_wl_r<104> a_wl_r<103> a_wl_r<102> a_wl_r<101> a_wl_r<100> a_wl_r<99> a_wl_r<98> a_wl_r<97> a_wl_r<96> a_wl_r<95> a_wl_r<94> a_wl_r<93> a_wl_r<92> a_wl_r<91> a_wl_r<90> a_wl_r<89> a_wl_r<88> a_wl_r<87> a_wl_r<86> a_wl_r<85> a_wl_r<84> a_wl_r<83> a_wl_r<82> a_wl_r<81> a_wl_r<80> a_wl_r<79> a_wl_r<78> a_wl_r<77> a_wl_r<76> a_wl_r<75> a_wl_r<74> a_wl_r<73> a_wl_r<72> a_wl_r<71> a_wl_r<70> a_wl_r<69> a_wl_r<68> a_wl_r<67> a_wl_r<66> a_wl_r<65> a_wl_r<64> a_wl_r<63> a_wl_r<62> a_wl_r<61> a_wl_r<60> a_wl_r<59> a_wl_r<58> a_wl_r<57> a_wl_r<56> a_wl_r<55> a_wl_r<54> a_wl_r<53> a_wl_r<52> a_wl_r<51> a_wl_r<50> a_wl_r<49> a_wl_r<48> a_wl_r<47> a_wl_r<46> a_wl_r<45> a_wl_r<44> a_wl_r<43> a_wl_r<42> a_wl_r<41> a_wl_r<40> a_wl_r<39> a_wl_r<38> a_wl_r<37> a_wl_r<36> a_wl_r<35> a_wl_r<34> a_wl_r<33> a_wl_r<32> a_wl_r<31> a_wl_r<30> a_wl_r<29> a_wl_r<28> a_wl_r<27> a_wl_r<26> a_wl_r<25> a_wl_r<24> a_wl_r<23> a_wl_r<22> a_wl_r<21> a_wl_r<20> a_wl_r<19> a_wl_r<18> a_wl_r<17> a_wl_r<16> a_wl_r<15> a_wl_r<14> a_wl_r<13> a_wl_r<12> a_wl_r<11> a_wl_r<10> a_wl_r<9> a_wl_r<8> a_wl_r<7> a_wl_r<6> a_wl_r<5> a_wl_r<4> a_wl_r<3> a_wl_r<2> a_wl_r<1> a_wl_r<0> VDDARRAY! VSS! / RM_IHPSG13_1024x64_c2_1P_MATRIX_pcell_1
XRAM<0> a_blc_l<127> a_blc_l<126> a_blc_l<125> a_blc_l<124> a_blc_l<123> a_blc_l<122> a_blc_l<121> a_blc_l<120> a_blc_l<119> a_blc_l<118> a_blc_l<117> a_blc_l<116> a_blc_l<115> a_blc_l<114> a_blc_l<113> a_blc_l<112> a_blc_l<111> a_blc_l<110> a_blc_l<109> a_blc_l<108> a_blc_l<107> a_blc_l<106> a_blc_l<105> a_blc_l<104> a_blc_l<103> a_blc_l<102> a_blc_l<101> a_blc_l<100> a_blc_l<99> a_blc_l<98> a_blc_l<97> a_blc_l<96> a_blc_l<95> a_blc_l<94> a_blc_l<93> a_blc_l<92> a_blc_l<91> a_blc_l<90> a_blc_l<89> a_blc_l<88> a_blc_l<87> a_blc_l<86> a_blc_l<85> a_blc_l<84> a_blc_l<83> a_blc_l<82> a_blc_l<81> a_blc_l<80> a_blc_l<79> a_blc_l<78> a_blc_l<77> a_blc_l<76> a_blc_l<75> a_blc_l<74> a_blc_l<73> a_blc_l<72> a_blc_l<71> a_blc_l<70> a_blc_l<69> a_blc_l<68> a_blc_l<67> a_blc_l<66> a_blc_l<65> a_blc_l<64> a_blc_l<63> a_blc_l<62> a_blc_l<61> a_blc_l<60> a_blc_l<59> a_blc_l<58> a_blc_l<57> a_blc_l<56> a_blc_l<55> a_blc_l<54> a_blc_l<53> a_blc_l<52> a_blc_l<51> a_blc_l<50> a_blc_l<49> a_blc_l<48> a_blc_l<47> a_blc_l<46> a_blc_l<45> a_blc_l<44> a_blc_l<43> a_blc_l<42> a_blc_l<41> a_blc_l<40> a_blc_l<39> a_blc_l<38> a_blc_l<37> a_blc_l<36> a_blc_l<35> a_blc_l<34> a_blc_l<33> a_blc_l<32> a_blc_l<31> a_blc_l<30> a_blc_l<29> a_blc_l<28> a_blc_l<27> a_blc_l<26> a_blc_l<25> a_blc_l<24> a_blc_l<23> a_blc_l<22> a_blc_l<21> a_blc_l<20> a_blc_l<19> a_blc_l<18> a_blc_l<17> a_blc_l<16> a_blc_l<15> a_blc_l<14> a_blc_l<13> a_blc_l<12> a_blc_l<11> a_blc_l<10> a_blc_l<9> a_blc_l<8> a_blc_l<7> a_blc_l<6> a_blc_l<5> a_blc_l<4> a_blc_l<3> a_blc_l<2> a_blc_l<1> a_blc_l<0> a_blt_l<127> a_blt_l<126> a_blt_l<125> a_blt_l<124> a_blt_l<123> a_blt_l<122> a_blt_l<121> a_blt_l<120> a_blt_l<119> a_blt_l<118> a_blt_l<117> a_blt_l<116> a_blt_l<115> a_blt_l<114> a_blt_l<113> a_blt_l<112> a_blt_l<111> a_blt_l<110> a_blt_l<109> a_blt_l<108> a_blt_l<107> a_blt_l<106> a_blt_l<105> a_blt_l<104> a_blt_l<103> a_blt_l<102> a_blt_l<101> a_blt_l<100> a_blt_l<99> a_blt_l<98> a_blt_l<97> a_blt_l<96> a_blt_l<95> a_blt_l<94> a_blt_l<93> a_blt_l<92> a_blt_l<91> a_blt_l<90> a_blt_l<89> a_blt_l<88> a_blt_l<87> a_blt_l<86> a_blt_l<85> a_blt_l<84> a_blt_l<83> a_blt_l<82> a_blt_l<81> a_blt_l<80> a_blt_l<79> a_blt_l<78> a_blt_l<77> a_blt_l<76> a_blt_l<75> a_blt_l<74> a_blt_l<73> a_blt_l<72> a_blt_l<71> a_blt_l<70> a_blt_l<69> a_blt_l<68> a_blt_l<67> a_blt_l<66> a_blt_l<65> a_blt_l<64> a_blt_l<63> a_blt_l<62> a_blt_l<61> a_blt_l<60> a_blt_l<59> a_blt_l<58> a_blt_l<57> a_blt_l<56> a_blt_l<55> a_blt_l<54> a_blt_l<53> a_blt_l<52> a_blt_l<51> a_blt_l<50> a_blt_l<49> a_blt_l<48> a_blt_l<47> a_blt_l<46> a_blt_l<45> a_blt_l<44> a_blt_l<43> a_blt_l<42> a_blt_l<41> a_blt_l<40> a_blt_l<39> a_blt_l<38> a_blt_l<37> a_blt_l<36> a_blt_l<35> a_blt_l<34> a_blt_l<33> a_blt_l<32> a_blt_l<31> a_blt_l<30> a_blt_l<29> a_blt_l<28> a_blt_l<27> a_blt_l<26> a_blt_l<25> a_blt_l<24> a_blt_l<23> a_blt_l<22> a_blt_l<21> a_blt_l<20> a_blt_l<19> a_blt_l<18> a_blt_l<17> a_blt_l<16> a_blt_l<15> a_blt_l<14> a_blt_l<13> a_blt_l<12> a_blt_l<11> a_blt_l<10> a_blt_l<9> a_blt_l<8> a_blt_l<7> a_blt_l<6> a_blt_l<5> a_blt_l<4> a_blt_l<3> a_blt_l<2> a_blt_l<1> a_blt_l<0> a_wl_l<255> a_wl_l<254> a_wl_l<253> a_wl_l<252> a_wl_l<251> a_wl_l<250> a_wl_l<249> a_wl_l<248> a_wl_l<247> a_wl_l<246> a_wl_l<245> a_wl_l<244> a_wl_l<243> a_wl_l<242> a_wl_l<241> a_wl_l<240> a_wl_l<239> a_wl_l<238> a_wl_l<237> a_wl_l<236> a_wl_l<235> a_wl_l<234> a_wl_l<233> a_wl_l<232> a_wl_l<231> a_wl_l<230> a_wl_l<229> a_wl_l<228> a_wl_l<227> a_wl_l<226> a_wl_l<225> a_wl_l<224> a_wl_l<223> a_wl_l<222> a_wl_l<221> a_wl_l<220> a_wl_l<219> a_wl_l<218> a_wl_l<217> a_wl_l<216> a_wl_l<215> a_wl_l<214> a_wl_l<213> a_wl_l<212> a_wl_l<211> a_wl_l<210> a_wl_l<209> a_wl_l<208> a_wl_l<207> a_wl_l<206> a_wl_l<205> a_wl_l<204> a_wl_l<203> a_wl_l<202> a_wl_l<201> a_wl_l<200> a_wl_l<199> a_wl_l<198> a_wl_l<197> a_wl_l<196> a_wl_l<195> a_wl_l<194> a_wl_l<193> a_wl_l<192> a_wl_l<191> a_wl_l<190> a_wl_l<189> a_wl_l<188> a_wl_l<187> a_wl_l<186> a_wl_l<185> a_wl_l<184> a_wl_l<183> a_wl_l<182> a_wl_l<181> a_wl_l<180> a_wl_l<179> a_wl_l<178> a_wl_l<177> a_wl_l<176> a_wl_l<175> a_wl_l<174> a_wl_l<173> a_wl_l<172> a_wl_l<171> a_wl_l<170> a_wl_l<169> a_wl_l<168> a_wl_l<167> a_wl_l<166> a_wl_l<165> a_wl_l<164> a_wl_l<163> a_wl_l<162> a_wl_l<161> a_wl_l<160> a_wl_l<159> a_wl_l<158> a_wl_l<157> a_wl_l<156> a_wl_l<155> a_wl_l<154> a_wl_l<153> a_wl_l<152> a_wl_l<151> a_wl_l<150> a_wl_l<149> a_wl_l<148> a_wl_l<147> a_wl_l<146> a_wl_l<145> a_wl_l<144> a_wl_l<143> a_wl_l<142> a_wl_l<141> a_wl_l<140> a_wl_l<139> a_wl_l<138> a_wl_l<137> a_wl_l<136> a_wl_l<135> a_wl_l<134> a_wl_l<133> a_wl_l<132> a_wl_l<131> a_wl_l<130> a_wl_l<129> a_wl_l<128> a_wl_l<127> a_wl_l<126> a_wl_l<125> a_wl_l<124> a_wl_l<123> a_wl_l<122> a_wl_l<121> a_wl_l<120> a_wl_l<119> a_wl_l<118> a_wl_l<117> a_wl_l<116> a_wl_l<115> a_wl_l<114> a_wl_l<113> a_wl_l<112> a_wl_l<111> a_wl_l<110> a_wl_l<109> a_wl_l<108> a_wl_l<107> a_wl_l<106> a_wl_l<105> a_wl_l<104> a_wl_l<103> a_wl_l<102> a_wl_l<101> a_wl_l<100> a_wl_l<99> a_wl_l<98> a_wl_l<97> a_wl_l<96> a_wl_l<95> a_wl_l<94> a_wl_l<93> a_wl_l<92> a_wl_l<91> a_wl_l<90> a_wl_l<89> a_wl_l<88> a_wl_l<87> a_wl_l<86> a_wl_l<85> a_wl_l<84> a_wl_l<83> a_wl_l<82> a_wl_l<81> a_wl_l<80> a_wl_l<79> a_wl_l<78> a_wl_l<77> a_wl_l<76> a_wl_l<75> a_wl_l<74> a_wl_l<73> a_wl_l<72> a_wl_l<71> a_wl_l<70> a_wl_l<69> a_wl_l<68> a_wl_l<67> a_wl_l<66> a_wl_l<65> a_wl_l<64> a_wl_l<63> a_wl_l<62> a_wl_l<61> a_wl_l<60> a_wl_l<59> a_wl_l<58> a_wl_l<57> a_wl_l<56> a_wl_l<55> a_wl_l<54> a_wl_l<53> a_wl_l<52> a_wl_l<51> a_wl_l<50> a_wl_l<49> a_wl_l<48> a_wl_l<47> a_wl_l<46> a_wl_l<45> a_wl_l<44> a_wl_l<43> a_wl_l<42> a_wl_l<41> a_wl_l<40> a_wl_l<39> a_wl_l<38> a_wl_l<37> a_wl_l<36> a_wl_l<35> a_wl_l<34> a_wl_l<33> a_wl_l<32> a_wl_l<31> a_wl_l<30> a_wl_l<29> a_wl_l<28> a_wl_l<27> a_wl_l<26> a_wl_l<25> a_wl_l<24> a_wl_l<23> a_wl_l<22> a_wl_l<21> a_wl_l<20> a_wl_l<19> a_wl_l<18> a_wl_l<17> a_wl_l<16> a_wl_l<15> a_wl_l<14> a_wl_l<13> a_wl_l<12> a_wl_l<11> a_wl_l<10> a_wl_l<9> a_wl_l<8> a_wl_l<7> a_wl_l<6> a_wl_l<5> a_wl_l<4> a_wl_l<3> a_wl_l<2> a_wl_l<1> a_wl_l<0> VDDARRAY! VSS! / RM_IHPSG13_1024x64_c2_1P_MATRIX_pcell_1


XA_COLDRV<1> a_addr_col<1> a_addr_col<0> a_addr_col_r<1> a_addr_col_r<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> a_addr_dec_r<7> a_addr_dec_r<6> a_addr_dec_r<5> a_addr_dec_r<4> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> a_dclk a_dclk_p_r<0> a_rclk a_rclk_p_r<0> a_wclk a_wclk_p_r<0> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13X8
XA_COLDRV<0> a_addr_col<1> a_addr_col<0> a_addr_col_l<1> a_addr_col_l<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> a_addr_dec_l<7> a_addr_dec_l<6> a_addr_dec_l<5> a_addr_dec_l<4> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> a_dclk a_dclk_p_l<0> a_rclk a_rclk_p_l<0> a_wclk a_wclk_p_l<0> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13X8


XA_WLDRV<31> a_wi<255> a_wi<254> a_wi<253> a_wi<252> a_wi<251> a_wi<250> a_wi<249> a_wi<248> a_wi<247> a_wi<246> a_wi<245> a_wi<244> a_wi<243> a_wi<242> a_wi<241> a_wi<240> a_wl_r<255> a_wl_r<254> a_wl_r<253> a_wl_r<252> a_wl_r<251> a_wl_r<250> a_wl_r<249> a_wl_r<248> a_wl_r<247> a_wl_r<246> a_wl_r<245> a_wl_r<244> a_wl_r<243> a_wl_r<242> a_wl_r<241> a_wl_r<240>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<30> a_wi<239> a_wi<238> a_wi<237> a_wi<236> a_wi<235> a_wi<234> a_wi<233> a_wi<232> a_wi<231> a_wi<230> a_wi<229> a_wi<228> a_wi<227> a_wi<226> a_wi<225> a_wi<224> a_wl_r<239> a_wl_r<238> a_wl_r<237> a_wl_r<236> a_wl_r<235> a_wl_r<234> a_wl_r<233> a_wl_r<232> a_wl_r<231> a_wl_r<230> a_wl_r<229> a_wl_r<228> a_wl_r<227> a_wl_r<226> a_wl_r<225> a_wl_r<224>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<29> a_wi<223> a_wi<222> a_wi<221> a_wi<220> a_wi<219> a_wi<218> a_wi<217> a_wi<216> a_wi<215> a_wi<214> a_wi<213> a_wi<212> a_wi<211> a_wi<210> a_wi<209> a_wi<208> a_wl_r<223> a_wl_r<222> a_wl_r<221> a_wl_r<220> a_wl_r<219> a_wl_r<218> a_wl_r<217> a_wl_r<216> a_wl_r<215> a_wl_r<214> a_wl_r<213> a_wl_r<212> a_wl_r<211> a_wl_r<210> a_wl_r<209> a_wl_r<208>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<28> a_wi<207> a_wi<206> a_wi<205> a_wi<204> a_wi<203> a_wi<202> a_wi<201> a_wi<200> a_wi<199> a_wi<198> a_wi<197> a_wi<196> a_wi<195> a_wi<194> a_wi<193> a_wi<192> a_wl_r<207> a_wl_r<206> a_wl_r<205> a_wl_r<204> a_wl_r<203> a_wl_r<202> a_wl_r<201> a_wl_r<200> a_wl_r<199> a_wl_r<198> a_wl_r<197> a_wl_r<196> a_wl_r<195> a_wl_r<194> a_wl_r<193> a_wl_r<192>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<27> a_wi<191> a_wi<190> a_wi<189> a_wi<188> a_wi<187> a_wi<186> a_wi<185> a_wi<184> a_wi<183> a_wi<182> a_wi<181> a_wi<180> a_wi<179> a_wi<178> a_wi<177> a_wi<176> a_wl_r<191> a_wl_r<190> a_wl_r<189> a_wl_r<188> a_wl_r<187> a_wl_r<186> a_wl_r<185> a_wl_r<184> a_wl_r<183> a_wl_r<182> a_wl_r<181> a_wl_r<180> a_wl_r<179> a_wl_r<178> a_wl_r<177> a_wl_r<176>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<26> a_wi<175> a_wi<174> a_wi<173> a_wi<172> a_wi<171> a_wi<170> a_wi<169> a_wi<168> a_wi<167> a_wi<166> a_wi<165> a_wi<164> a_wi<163> a_wi<162> a_wi<161> a_wi<160> a_wl_r<175> a_wl_r<174> a_wl_r<173> a_wl_r<172> a_wl_r<171> a_wl_r<170> a_wl_r<169> a_wl_r<168> a_wl_r<167> a_wl_r<166> a_wl_r<165> a_wl_r<164> a_wl_r<163> a_wl_r<162> a_wl_r<161> a_wl_r<160>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<25> a_wi<159> a_wi<158> a_wi<157> a_wi<156> a_wi<155> a_wi<154> a_wi<153> a_wi<152> a_wi<151> a_wi<150> a_wi<149> a_wi<148> a_wi<147> a_wi<146> a_wi<145> a_wi<144> a_wl_r<159> a_wl_r<158> a_wl_r<157> a_wl_r<156> a_wl_r<155> a_wl_r<154> a_wl_r<153> a_wl_r<152> a_wl_r<151> a_wl_r<150> a_wl_r<149> a_wl_r<148> a_wl_r<147> a_wl_r<146> a_wl_r<145> a_wl_r<144>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<24> a_wi<143> a_wi<142> a_wi<141> a_wi<140> a_wi<139> a_wi<138> a_wi<137> a_wi<136> a_wi<135> a_wi<134> a_wi<133> a_wi<132> a_wi<131> a_wi<130> a_wi<129> a_wi<128> a_wl_r<143> a_wl_r<142> a_wl_r<141> a_wl_r<140> a_wl_r<139> a_wl_r<138> a_wl_r<137> a_wl_r<136> a_wl_r<135> a_wl_r<134> a_wl_r<133> a_wl_r<132> a_wl_r<131> a_wl_r<130> a_wl_r<129> a_wl_r<128>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<23> a_wi<127> a_wi<126> a_wi<125> a_wi<124> a_wi<123> a_wi<122> a_wi<121> a_wi<120> a_wi<119> a_wi<118> a_wi<117> a_wi<116> a_wi<115> a_wi<114> a_wi<113> a_wi<112> a_wl_r<127> a_wl_r<126> a_wl_r<125> a_wl_r<124> a_wl_r<123> a_wl_r<122> a_wl_r<121> a_wl_r<120> a_wl_r<119> a_wl_r<118> a_wl_r<117> a_wl_r<116> a_wl_r<115> a_wl_r<114> a_wl_r<113> a_wl_r<112>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<22> a_wi<111> a_wi<110> a_wi<109> a_wi<108> a_wi<107> a_wi<106> a_wi<105> a_wi<104> a_wi<103> a_wi<102> a_wi<101> a_wi<100> a_wi<99> a_wi<98> a_wi<97> a_wi<96> a_wl_r<111> a_wl_r<110> a_wl_r<109> a_wl_r<108> a_wl_r<107> a_wl_r<106> a_wl_r<105> a_wl_r<104> a_wl_r<103> a_wl_r<102> a_wl_r<101> a_wl_r<100> a_wl_r<99> a_wl_r<98> a_wl_r<97> a_wl_r<96>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<21> a_wi<95> a_wi<94> a_wi<93> a_wi<92> a_wi<91> a_wi<90> a_wi<89> a_wi<88> a_wi<87> a_wi<86> a_wi<85> a_wi<84> a_wi<83> a_wi<82> a_wi<81> a_wi<80> a_wl_r<95> a_wl_r<94> a_wl_r<93> a_wl_r<92> a_wl_r<91> a_wl_r<90> a_wl_r<89> a_wl_r<88> a_wl_r<87> a_wl_r<86> a_wl_r<85> a_wl_r<84> a_wl_r<83> a_wl_r<82> a_wl_r<81> a_wl_r<80>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<20> a_wi<79> a_wi<78> a_wi<77> a_wi<76> a_wi<75> a_wi<74> a_wi<73> a_wi<72> a_wi<71> a_wi<70> a_wi<69> a_wi<68> a_wi<67> a_wi<66> a_wi<65> a_wi<64> a_wl_r<79> a_wl_r<78> a_wl_r<77> a_wl_r<76> a_wl_r<75> a_wl_r<74> a_wl_r<73> a_wl_r<72> a_wl_r<71> a_wl_r<70> a_wl_r<69> a_wl_r<68> a_wl_r<67> a_wl_r<66> a_wl_r<65> a_wl_r<64>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<19> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wl_r<63> a_wl_r<62> a_wl_r<61> a_wl_r<60> a_wl_r<59> a_wl_r<58> a_wl_r<57> a_wl_r<56> a_wl_r<55> a_wl_r<54> a_wl_r<53> a_wl_r<52> a_wl_r<51> a_wl_r<50> a_wl_r<49> a_wl_r<48>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<18> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wl_r<47> a_wl_r<46> a_wl_r<45> a_wl_r<44> a_wl_r<43> a_wl_r<42> a_wl_r<41> a_wl_r<40> a_wl_r<39> a_wl_r<38> a_wl_r<37> a_wl_r<36> a_wl_r<35> a_wl_r<34> a_wl_r<33> a_wl_r<32>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<17> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wl_r<31> a_wl_r<30> a_wl_r<29> a_wl_r<28> a_wl_r<27> a_wl_r<26> a_wl_r<25> a_wl_r<24> a_wl_r<23> a_wl_r<22> a_wl_r<21> a_wl_r<20> a_wl_r<19> a_wl_r<18> a_wl_r<17> a_wl_r<16>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<16> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> a_wl_r<15> a_wl_r<14> a_wl_r<13> a_wl_r<12> a_wl_r<11> a_wl_r<10> a_wl_r<9> a_wl_r<8> a_wl_r<7> a_wl_r<6> a_wl_r<5> a_wl_r<4> a_wl_r<3> a_wl_r<2> a_wl_r<1> a_wl_r<0>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<15> a_wi<255> a_wi<254> a_wi<253> a_wi<252> a_wi<251> a_wi<250> a_wi<249> a_wi<248> a_wi<247> a_wi<246> a_wi<245> a_wi<244> a_wi<243> a_wi<242> a_wi<241> a_wi<240> a_wl_l<255> a_wl_l<254> a_wl_l<253> a_wl_l<252> a_wl_l<251> a_wl_l<250> a_wl_l<249> a_wl_l<248> a_wl_l<247> a_wl_l<246> a_wl_l<245> a_wl_l<244> a_wl_l<243> a_wl_l<242> a_wl_l<241> a_wl_l<240>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<14> a_wi<239> a_wi<238> a_wi<237> a_wi<236> a_wi<235> a_wi<234> a_wi<233> a_wi<232> a_wi<231> a_wi<230> a_wi<229> a_wi<228> a_wi<227> a_wi<226> a_wi<225> a_wi<224> a_wl_l<239> a_wl_l<238> a_wl_l<237> a_wl_l<236> a_wl_l<235> a_wl_l<234> a_wl_l<233> a_wl_l<232> a_wl_l<231> a_wl_l<230> a_wl_l<229> a_wl_l<228> a_wl_l<227> a_wl_l<226> a_wl_l<225> a_wl_l<224>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<13> a_wi<223> a_wi<222> a_wi<221> a_wi<220> a_wi<219> a_wi<218> a_wi<217> a_wi<216> a_wi<215> a_wi<214> a_wi<213> a_wi<212> a_wi<211> a_wi<210> a_wi<209> a_wi<208> a_wl_l<223> a_wl_l<222> a_wl_l<221> a_wl_l<220> a_wl_l<219> a_wl_l<218> a_wl_l<217> a_wl_l<216> a_wl_l<215> a_wl_l<214> a_wl_l<213> a_wl_l<212> a_wl_l<211> a_wl_l<210> a_wl_l<209> a_wl_l<208>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<12> a_wi<207> a_wi<206> a_wi<205> a_wi<204> a_wi<203> a_wi<202> a_wi<201> a_wi<200> a_wi<199> a_wi<198> a_wi<197> a_wi<196> a_wi<195> a_wi<194> a_wi<193> a_wi<192> a_wl_l<207> a_wl_l<206> a_wl_l<205> a_wl_l<204> a_wl_l<203> a_wl_l<202> a_wl_l<201> a_wl_l<200> a_wl_l<199> a_wl_l<198> a_wl_l<197> a_wl_l<196> a_wl_l<195> a_wl_l<194> a_wl_l<193> a_wl_l<192>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<11> a_wi<191> a_wi<190> a_wi<189> a_wi<188> a_wi<187> a_wi<186> a_wi<185> a_wi<184> a_wi<183> a_wi<182> a_wi<181> a_wi<180> a_wi<179> a_wi<178> a_wi<177> a_wi<176> a_wl_l<191> a_wl_l<190> a_wl_l<189> a_wl_l<188> a_wl_l<187> a_wl_l<186> a_wl_l<185> a_wl_l<184> a_wl_l<183> a_wl_l<182> a_wl_l<181> a_wl_l<180> a_wl_l<179> a_wl_l<178> a_wl_l<177> a_wl_l<176>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<10> a_wi<175> a_wi<174> a_wi<173> a_wi<172> a_wi<171> a_wi<170> a_wi<169> a_wi<168> a_wi<167> a_wi<166> a_wi<165> a_wi<164> a_wi<163> a_wi<162> a_wi<161> a_wi<160> a_wl_l<175> a_wl_l<174> a_wl_l<173> a_wl_l<172> a_wl_l<171> a_wl_l<170> a_wl_l<169> a_wl_l<168> a_wl_l<167> a_wl_l<166> a_wl_l<165> a_wl_l<164> a_wl_l<163> a_wl_l<162> a_wl_l<161> a_wl_l<160>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<9> a_wi<159> a_wi<158> a_wi<157> a_wi<156> a_wi<155> a_wi<154> a_wi<153> a_wi<152> a_wi<151> a_wi<150> a_wi<149> a_wi<148> a_wi<147> a_wi<146> a_wi<145> a_wi<144> a_wl_l<159> a_wl_l<158> a_wl_l<157> a_wl_l<156> a_wl_l<155> a_wl_l<154> a_wl_l<153> a_wl_l<152> a_wl_l<151> a_wl_l<150> a_wl_l<149> a_wl_l<148> a_wl_l<147> a_wl_l<146> a_wl_l<145> a_wl_l<144>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<8> a_wi<143> a_wi<142> a_wi<141> a_wi<140> a_wi<139> a_wi<138> a_wi<137> a_wi<136> a_wi<135> a_wi<134> a_wi<133> a_wi<132> a_wi<131> a_wi<130> a_wi<129> a_wi<128> a_wl_l<143> a_wl_l<142> a_wl_l<141> a_wl_l<140> a_wl_l<139> a_wl_l<138> a_wl_l<137> a_wl_l<136> a_wl_l<135> a_wl_l<134> a_wl_l<133> a_wl_l<132> a_wl_l<131> a_wl_l<130> a_wl_l<129> a_wl_l<128>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<7> a_wi<127> a_wi<126> a_wi<125> a_wi<124> a_wi<123> a_wi<122> a_wi<121> a_wi<120> a_wi<119> a_wi<118> a_wi<117> a_wi<116> a_wi<115> a_wi<114> a_wi<113> a_wi<112> a_wl_l<127> a_wl_l<126> a_wl_l<125> a_wl_l<124> a_wl_l<123> a_wl_l<122> a_wl_l<121> a_wl_l<120> a_wl_l<119> a_wl_l<118> a_wl_l<117> a_wl_l<116> a_wl_l<115> a_wl_l<114> a_wl_l<113> a_wl_l<112>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<6> a_wi<111> a_wi<110> a_wi<109> a_wi<108> a_wi<107> a_wi<106> a_wi<105> a_wi<104> a_wi<103> a_wi<102> a_wi<101> a_wi<100> a_wi<99> a_wi<98> a_wi<97> a_wi<96> a_wl_l<111> a_wl_l<110> a_wl_l<109> a_wl_l<108> a_wl_l<107> a_wl_l<106> a_wl_l<105> a_wl_l<104> a_wl_l<103> a_wl_l<102> a_wl_l<101> a_wl_l<100> a_wl_l<99> a_wl_l<98> a_wl_l<97> a_wl_l<96>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<5> a_wi<95> a_wi<94> a_wi<93> a_wi<92> a_wi<91> a_wi<90> a_wi<89> a_wi<88> a_wi<87> a_wi<86> a_wi<85> a_wi<84> a_wi<83> a_wi<82> a_wi<81> a_wi<80> a_wl_l<95> a_wl_l<94> a_wl_l<93> a_wl_l<92> a_wl_l<91> a_wl_l<90> a_wl_l<89> a_wl_l<88> a_wl_l<87> a_wl_l<86> a_wl_l<85> a_wl_l<84> a_wl_l<83> a_wl_l<82> a_wl_l<81> a_wl_l<80>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<4> a_wi<79> a_wi<78> a_wi<77> a_wi<76> a_wi<75> a_wi<74> a_wi<73> a_wi<72> a_wi<71> a_wi<70> a_wi<69> a_wi<68> a_wi<67> a_wi<66> a_wi<65> a_wi<64> a_wl_l<79> a_wl_l<78> a_wl_l<77> a_wl_l<76> a_wl_l<75> a_wl_l<74> a_wl_l<73> a_wl_l<72> a_wl_l<71> a_wl_l<70> a_wl_l<69> a_wl_l<68> a_wl_l<67> a_wl_l<66> a_wl_l<65> a_wl_l<64>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<3> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wl_l<63> a_wl_l<62> a_wl_l<61> a_wl_l<60> a_wl_l<59> a_wl_l<58> a_wl_l<57> a_wl_l<56> a_wl_l<55> a_wl_l<54> a_wl_l<53> a_wl_l<52> a_wl_l<51> a_wl_l<50> a_wl_l<49> a_wl_l<48>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<2> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wl_l<47> a_wl_l<46> a_wl_l<45> a_wl_l<44> a_wl_l<43> a_wl_l<42> a_wl_l<41> a_wl_l<40> a_wl_l<39> a_wl_l<38> a_wl_l<37> a_wl_l<36> a_wl_l<35> a_wl_l<34> a_wl_l<33> a_wl_l<32>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<1> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wl_l<31> a_wl_l<30> a_wl_l<29> a_wl_l<28> a_wl_l<27> a_wl_l<26> a_wl_l<25> a_wl_l<24> a_wl_l<23> a_wl_l<22> a_wl_l<21> a_wl_l<20> a_wl_l<19> a_wl_l<18> a_wl_l<17> a_wl_l<16>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8
XA_WLDRV<0> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> a_wl_l<15> a_wl_l<14> a_wl_l<13> a_wl_l<12> a_wl_l<11> a_wl_l<10> a_wl_l<9> a_wl_l<8> a_wl_l<7> a_wl_l<6> a_wl_l<5> a_wl_l<4> a_wl_l<3> a_wl_l<2> a_wl_l<1> a_wl_l<0>  VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_WLDRV16X8


XA_CTRL a_aclk_n A_BIST_CLK A_BIST_MEN A_BIST_EN A_BIST_REN A_BIST_WEN a_tiel A_CLK A_MEN a_dclk a_eclk a_pulse_h a_pulse_l a_pulse a_rclk A_REN a_cs a_wclk A_WEN VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_CTRL


XA_ROWDEC a_addr_row<7> a_addr_row<6> a_addr_row<5> a_addr_row<4> a_addr_row<3> a_addr_row<2> a_addr_row<1> a_addr_row<0> a_cs a_eclk a_wi<255> a_wi<254> a_wi<253> a_wi<252> a_wi<251> a_wi<250> a_wi<249> a_wi<248> a_wi<247> a_wi<246> a_wi<245> a_wi<244> a_wi<243> a_wi<242> a_wi<241> a_wi<240> a_wi<239> a_wi<238> a_wi<237> a_wi<236> a_wi<235> a_wi<234> a_wi<233> a_wi<232> a_wi<231> a_wi<230> a_wi<229> a_wi<228> a_wi<227> a_wi<226> a_wi<225> a_wi<224> a_wi<223> a_wi<222> a_wi<221> a_wi<220> a_wi<219> a_wi<218> a_wi<217> a_wi<216> a_wi<215> a_wi<214> a_wi<213> a_wi<212> a_wi<211> a_wi<210> a_wi<209> a_wi<208> a_wi<207> a_wi<206> a_wi<205> a_wi<204> a_wi<203> a_wi<202> a_wi<201> a_wi<200> a_wi<199> a_wi<198> a_wi<197> a_wi<196> a_wi<195> a_wi<194> a_wi<193> a_wi<192> a_wi<191> a_wi<190> a_wi<189> a_wi<188> a_wi<187> a_wi<186> a_wi<185> a_wi<184> a_wi<183> a_wi<182> a_wi<181> a_wi<180> a_wi<179> a_wi<178> a_wi<177> a_wi<176> a_wi<175> a_wi<174> a_wi<173> a_wi<172> a_wi<171> a_wi<170> a_wi<169> a_wi<168> a_wi<167> a_wi<166> a_wi<165> a_wi<164> a_wi<163> a_wi<162> a_wi<161> a_wi<160> a_wi<159> a_wi<158> a_wi<157> a_wi<156> a_wi<155> a_wi<154> a_wi<153> a_wi<152> a_wi<151> a_wi<150> a_wi<149> a_wi<148> a_wi<147> a_wi<146> a_wi<145> a_wi<144> a_wi<143> a_wi<142> a_wi<141> a_wi<140> a_wi<139> a_wi<138> a_wi<137> a_wi<136> a_wi<135> a_wi<134> a_wi<133> a_wi<132> a_wi<131> a_wi<130> a_wi<129> a_wi<128> a_wi<127> a_wi<126> a_wi<125> a_wi<124> a_wi<123> a_wi<122> a_wi<121> a_wi<120> a_wi<119> a_wi<118> a_wi<117> a_wi<116> a_wi<115> a_wi<114> a_wi<113> a_wi<112> a_wi<111> a_wi<110> a_wi<109> a_wi<108> a_wi<107> a_wi<106> a_wi<105> a_wi<104> a_wi<103> a_wi<102> a_wi<101> a_wi<100> a_wi<99> a_wi<98> a_wi<97> a_wi<96> a_wi<95> a_wi<94> a_wi<93> a_wi<92> a_wi<91> a_wi<90> a_wi<89> a_wi<88> a_wi<87> a_wi<86> a_wi<85> a_wi<84> a_wi<83> a_wi<82> a_wi<81> a_wi<80> a_wi<79> a_wi<78> a_wi<77> a_wi<76> a_wi<75> a_wi<74> a_wi<73> a_wi<72> a_wi<71> a_wi<70> a_wi<69> a_wi<68> a_wi<67> a_wi<66> a_wi<65> a_wi<64> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_ROWDEC8
XA_ROWREG a_aclk_n A_ADDR<9> A_ADDR<8> A_ADDR<7> A_ADDR<6> A_ADDR<5> A_ADDR<4> A_ADDR<3> A_ADDR<2> a_addr_row<7> a_addr_row<6> a_addr_row<5> a_addr_row<4> a_addr_row<3> a_addr_row<2> a_addr_row<1> a_addr_row<0> A_BIST_ADDR<9> A_BIST_ADDR<8> A_BIST_ADDR<7> A_BIST_ADDR<6> A_BIST_ADDR<5> A_BIST_ADDR<4> A_BIST_ADDR<3> A_BIST_ADDR<2> A_BIST_EN VDD! VSS!  / RM_IHPSG13_1024x64_c2_1P_ROWREG8
XA_COLDEC a_aclk_n A_ADDR<1> A_ADDR<0> a_addr_col<1> a_addr_col<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> A_BIST_ADDR<1> A_BIST_ADDR<0> A_BIST_EN VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDEC2


XA_DLYH a_pulse a_pulse_h VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_DLY_pcell_2
XA_DLYL a_pulse_x a_pulse_l VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_DLY_pcell_3
XA_DLYMUX a_pulse_h A_DLY a_pulse_x VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_DLY_MUX

XCOLCTRL<63> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<63> A_BIST_DIN<63> A_BIST_EN a_blc_r<127> a_blc_r<126> a_blc_r<125> a_blc_r<124> a_blt_r<127> a_blt_r<126> a_blt_r<125> a_blt_r<124> A_BM<63> a_dclk_n_r<31> a_dclk_n_r<32> a_dclk_p_r<31> a_dclk_p_r<32> A_DOUT<63> A_DIN<63> a_rclk_n_r<31> a_rclk_n_r<32> a_rclk_p_r<31> a_rclk_p_r<32> a_tieh<63> a_wclk_n_r<31> a_wclk_n_r<32> a_wclk_p_r<31> a_wclk_p_r<32> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<62> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<62> A_BIST_DIN<62> A_BIST_EN a_blc_r<123> a_blc_r<122> a_blc_r<121> a_blc_r<120> a_blt_r<123> a_blt_r<122> a_blt_r<121> a_blt_r<120> A_BM<62> a_dclk_n_r<30> a_dclk_n_r<31> a_dclk_p_r<30> a_dclk_p_r<31> A_DOUT<62> A_DIN<62> a_rclk_n_r<30> a_rclk_n_r<31> a_rclk_p_r<30> a_rclk_p_r<31> a_tieh<62> a_wclk_n_r<30> a_wclk_n_r<31> a_wclk_p_r<30> a_wclk_p_r<31> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<61> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<61> A_BIST_DIN<61> A_BIST_EN a_blc_r<119> a_blc_r<118> a_blc_r<117> a_blc_r<116> a_blt_r<119> a_blt_r<118> a_blt_r<117> a_blt_r<116> A_BM<61> a_dclk_n_r<29> a_dclk_n_r<30> a_dclk_p_r<29> a_dclk_p_r<30> A_DOUT<61> A_DIN<61> a_rclk_n_r<29> a_rclk_n_r<30> a_rclk_p_r<29> a_rclk_p_r<30> a_tieh<61> a_wclk_n_r<29> a_wclk_n_r<30> a_wclk_p_r<29> a_wclk_p_r<30> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<60> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<60> A_BIST_DIN<60> A_BIST_EN a_blc_r<115> a_blc_r<114> a_blc_r<113> a_blc_r<112> a_blt_r<115> a_blt_r<114> a_blt_r<113> a_blt_r<112> A_BM<60> a_dclk_n_r<28> a_dclk_n_r<29> a_dclk_p_r<28> a_dclk_p_r<29> A_DOUT<60> A_DIN<60> a_rclk_n_r<28> a_rclk_n_r<29> a_rclk_p_r<28> a_rclk_p_r<29> a_tieh<60> a_wclk_n_r<28> a_wclk_n_r<29> a_wclk_p_r<28> a_wclk_p_r<29> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<59> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<59> A_BIST_DIN<59> A_BIST_EN a_blc_r<111> a_blc_r<110> a_blc_r<109> a_blc_r<108> a_blt_r<111> a_blt_r<110> a_blt_r<109> a_blt_r<108> A_BM<59> a_dclk_n_r<27> a_dclk_n_r<28> a_dclk_p_r<27> a_dclk_p_r<28> A_DOUT<59> A_DIN<59> a_rclk_n_r<27> a_rclk_n_r<28> a_rclk_p_r<27> a_rclk_p_r<28> a_tieh<59> a_wclk_n_r<27> a_wclk_n_r<28> a_wclk_p_r<27> a_wclk_p_r<28> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<58> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<58> A_BIST_DIN<58> A_BIST_EN a_blc_r<107> a_blc_r<106> a_blc_r<105> a_blc_r<104> a_blt_r<107> a_blt_r<106> a_blt_r<105> a_blt_r<104> A_BM<58> a_dclk_n_r<26> a_dclk_n_r<27> a_dclk_p_r<26> a_dclk_p_r<27> A_DOUT<58> A_DIN<58> a_rclk_n_r<26> a_rclk_n_r<27> a_rclk_p_r<26> a_rclk_p_r<27> a_tieh<58> a_wclk_n_r<26> a_wclk_n_r<27> a_wclk_p_r<26> a_wclk_p_r<27> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<57> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<57> A_BIST_DIN<57> A_BIST_EN a_blc_r<103> a_blc_r<102> a_blc_r<101> a_blc_r<100> a_blt_r<103> a_blt_r<102> a_blt_r<101> a_blt_r<100> A_BM<57> a_dclk_n_r<25> a_dclk_n_r<26> a_dclk_p_r<25> a_dclk_p_r<26> A_DOUT<57> A_DIN<57> a_rclk_n_r<25> a_rclk_n_r<26> a_rclk_p_r<25> a_rclk_p_r<26> a_tieh<57> a_wclk_n_r<25> a_wclk_n_r<26> a_wclk_p_r<25> a_wclk_p_r<26> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<56> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<56> A_BIST_DIN<56> A_BIST_EN a_blc_r<99> a_blc_r<98> a_blc_r<97> a_blc_r<96> a_blt_r<99> a_blt_r<98> a_blt_r<97> a_blt_r<96> A_BM<56> a_dclk_n_r<24> a_dclk_n_r<25> a_dclk_p_r<24> a_dclk_p_r<25> A_DOUT<56> A_DIN<56> a_rclk_n_r<24> a_rclk_n_r<25> a_rclk_p_r<24> a_rclk_p_r<25> a_tieh<56> a_wclk_n_r<24> a_wclk_n_r<25> a_wclk_p_r<24> a_wclk_p_r<25> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<55> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<55> A_BIST_DIN<55> A_BIST_EN a_blc_r<95> a_blc_r<94> a_blc_r<93> a_blc_r<92> a_blt_r<95> a_blt_r<94> a_blt_r<93> a_blt_r<92> A_BM<55> a_dclk_n_r<23> a_dclk_n_r<24> a_dclk_p_r<23> a_dclk_p_r<24> A_DOUT<55> A_DIN<55> a_rclk_n_r<23> a_rclk_n_r<24> a_rclk_p_r<23> a_rclk_p_r<24> a_tieh<55> a_wclk_n_r<23> a_wclk_n_r<24> a_wclk_p_r<23> a_wclk_p_r<24> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<54> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<54> A_BIST_DIN<54> A_BIST_EN a_blc_r<91> a_blc_r<90> a_blc_r<89> a_blc_r<88> a_blt_r<91> a_blt_r<90> a_blt_r<89> a_blt_r<88> A_BM<54> a_dclk_n_r<22> a_dclk_n_r<23> a_dclk_p_r<22> a_dclk_p_r<23> A_DOUT<54> A_DIN<54> a_rclk_n_r<22> a_rclk_n_r<23> a_rclk_p_r<22> a_rclk_p_r<23> a_tieh<54> a_wclk_n_r<22> a_wclk_n_r<23> a_wclk_p_r<22> a_wclk_p_r<23> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<53> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<53> A_BIST_DIN<53> A_BIST_EN a_blc_r<87> a_blc_r<86> a_blc_r<85> a_blc_r<84> a_blt_r<87> a_blt_r<86> a_blt_r<85> a_blt_r<84> A_BM<53> a_dclk_n_r<21> a_dclk_n_r<22> a_dclk_p_r<21> a_dclk_p_r<22> A_DOUT<53> A_DIN<53> a_rclk_n_r<21> a_rclk_n_r<22> a_rclk_p_r<21> a_rclk_p_r<22> a_tieh<53> a_wclk_n_r<21> a_wclk_n_r<22> a_wclk_p_r<21> a_wclk_p_r<22> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<52> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<52> A_BIST_DIN<52> A_BIST_EN a_blc_r<83> a_blc_r<82> a_blc_r<81> a_blc_r<80> a_blt_r<83> a_blt_r<82> a_blt_r<81> a_blt_r<80> A_BM<52> a_dclk_n_r<20> a_dclk_n_r<21> a_dclk_p_r<20> a_dclk_p_r<21> A_DOUT<52> A_DIN<52> a_rclk_n_r<20> a_rclk_n_r<21> a_rclk_p_r<20> a_rclk_p_r<21> a_tieh<52> a_wclk_n_r<20> a_wclk_n_r<21> a_wclk_p_r<20> a_wclk_p_r<21> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<51> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<51> A_BIST_DIN<51> A_BIST_EN a_blc_r<79> a_blc_r<78> a_blc_r<77> a_blc_r<76> a_blt_r<79> a_blt_r<78> a_blt_r<77> a_blt_r<76> A_BM<51> a_dclk_n_r<19> a_dclk_n_r<20> a_dclk_p_r<19> a_dclk_p_r<20> A_DOUT<51> A_DIN<51> a_rclk_n_r<19> a_rclk_n_r<20> a_rclk_p_r<19> a_rclk_p_r<20> a_tieh<51> a_wclk_n_r<19> a_wclk_n_r<20> a_wclk_p_r<19> a_wclk_p_r<20> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<50> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<50> A_BIST_DIN<50> A_BIST_EN a_blc_r<75> a_blc_r<74> a_blc_r<73> a_blc_r<72> a_blt_r<75> a_blt_r<74> a_blt_r<73> a_blt_r<72> A_BM<50> a_dclk_n_r<18> a_dclk_n_r<19> a_dclk_p_r<18> a_dclk_p_r<19> A_DOUT<50> A_DIN<50> a_rclk_n_r<18> a_rclk_n_r<19> a_rclk_p_r<18> a_rclk_p_r<19> a_tieh<50> a_wclk_n_r<18> a_wclk_n_r<19> a_wclk_p_r<18> a_wclk_p_r<19> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<49> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<49> A_BIST_DIN<49> A_BIST_EN a_blc_r<71> a_blc_r<70> a_blc_r<69> a_blc_r<68> a_blt_r<71> a_blt_r<70> a_blt_r<69> a_blt_r<68> A_BM<49> a_dclk_n_r<17> a_dclk_n_r<18> a_dclk_p_r<17> a_dclk_p_r<18> A_DOUT<49> A_DIN<49> a_rclk_n_r<17> a_rclk_n_r<18> a_rclk_p_r<17> a_rclk_p_r<18> a_tieh<49> a_wclk_n_r<17> a_wclk_n_r<18> a_wclk_p_r<17> a_wclk_p_r<18> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<48> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<48> A_BIST_DIN<48> A_BIST_EN a_blc_r<67> a_blc_r<66> a_blc_r<65> a_blc_r<64> a_blt_r<67> a_blt_r<66> a_blt_r<65> a_blt_r<64> A_BM<48> a_dclk_n_r<16> a_dclk_n_r<17> a_dclk_p_r<16> a_dclk_p_r<17> A_DOUT<48> A_DIN<48> a_rclk_n_r<16> a_rclk_n_r<17> a_rclk_p_r<16> a_rclk_p_r<17> a_tieh<48> a_wclk_n_r<16> a_wclk_n_r<17> a_wclk_p_r<16> a_wclk_p_r<17> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<47> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<47> A_BIST_DIN<47> A_BIST_EN a_blc_r<63> a_blc_r<62> a_blc_r<61> a_blc_r<60> a_blt_r<63> a_blt_r<62> a_blt_r<61> a_blt_r<60> A_BM<47> a_dclk_n_r<15> a_dclk_n_r<16> a_dclk_p_r<15> a_dclk_p_r<16> A_DOUT<47> A_DIN<47> a_rclk_n_r<15> a_rclk_n_r<16> a_rclk_p_r<15> a_rclk_p_r<16> a_tieh<47> a_wclk_n_r<15> a_wclk_n_r<16> a_wclk_p_r<15> a_wclk_p_r<16> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<46> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<46> A_BIST_DIN<46> A_BIST_EN a_blc_r<59> a_blc_r<58> a_blc_r<57> a_blc_r<56> a_blt_r<59> a_blt_r<58> a_blt_r<57> a_blt_r<56> A_BM<46> a_dclk_n_r<14> a_dclk_n_r<15> a_dclk_p_r<14> a_dclk_p_r<15> A_DOUT<46> A_DIN<46> a_rclk_n_r<14> a_rclk_n_r<15> a_rclk_p_r<14> a_rclk_p_r<15> a_tieh<46> a_wclk_n_r<14> a_wclk_n_r<15> a_wclk_p_r<14> a_wclk_p_r<15> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<45> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<45> A_BIST_DIN<45> A_BIST_EN a_blc_r<55> a_blc_r<54> a_blc_r<53> a_blc_r<52> a_blt_r<55> a_blt_r<54> a_blt_r<53> a_blt_r<52> A_BM<45> a_dclk_n_r<13> a_dclk_n_r<14> a_dclk_p_r<13> a_dclk_p_r<14> A_DOUT<45> A_DIN<45> a_rclk_n_r<13> a_rclk_n_r<14> a_rclk_p_r<13> a_rclk_p_r<14> a_tieh<45> a_wclk_n_r<13> a_wclk_n_r<14> a_wclk_p_r<13> a_wclk_p_r<14> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<44> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<44> A_BIST_DIN<44> A_BIST_EN a_blc_r<51> a_blc_r<50> a_blc_r<49> a_blc_r<48> a_blt_r<51> a_blt_r<50> a_blt_r<49> a_blt_r<48> A_BM<44> a_dclk_n_r<12> a_dclk_n_r<13> a_dclk_p_r<12> a_dclk_p_r<13> A_DOUT<44> A_DIN<44> a_rclk_n_r<12> a_rclk_n_r<13> a_rclk_p_r<12> a_rclk_p_r<13> a_tieh<44> a_wclk_n_r<12> a_wclk_n_r<13> a_wclk_p_r<12> a_wclk_p_r<13> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<43> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<43> A_BIST_DIN<43> A_BIST_EN a_blc_r<47> a_blc_r<46> a_blc_r<45> a_blc_r<44> a_blt_r<47> a_blt_r<46> a_blt_r<45> a_blt_r<44> A_BM<43> a_dclk_n_r<11> a_dclk_n_r<12> a_dclk_p_r<11> a_dclk_p_r<12> A_DOUT<43> A_DIN<43> a_rclk_n_r<11> a_rclk_n_r<12> a_rclk_p_r<11> a_rclk_p_r<12> a_tieh<43> a_wclk_n_r<11> a_wclk_n_r<12> a_wclk_p_r<11> a_wclk_p_r<12> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<42> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<42> A_BIST_DIN<42> A_BIST_EN a_blc_r<43> a_blc_r<42> a_blc_r<41> a_blc_r<40> a_blt_r<43> a_blt_r<42> a_blt_r<41> a_blt_r<40> A_BM<42> a_dclk_n_r<10> a_dclk_n_r<11> a_dclk_p_r<10> a_dclk_p_r<11> A_DOUT<42> A_DIN<42> a_rclk_n_r<10> a_rclk_n_r<11> a_rclk_p_r<10> a_rclk_p_r<11> a_tieh<42> a_wclk_n_r<10> a_wclk_n_r<11> a_wclk_p_r<10> a_wclk_p_r<11> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<41> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<41> A_BIST_DIN<41> A_BIST_EN a_blc_r<39> a_blc_r<38> a_blc_r<37> a_blc_r<36> a_blt_r<39> a_blt_r<38> a_blt_r<37> a_blt_r<36> A_BM<41> a_dclk_n_r<9> a_dclk_n_r<10> a_dclk_p_r<9> a_dclk_p_r<10> A_DOUT<41> A_DIN<41> a_rclk_n_r<9> a_rclk_n_r<10> a_rclk_p_r<9> a_rclk_p_r<10> a_tieh<41> a_wclk_n_r<9> a_wclk_n_r<10> a_wclk_p_r<9> a_wclk_p_r<10> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<40> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<40> A_BIST_DIN<40> A_BIST_EN a_blc_r<35> a_blc_r<34> a_blc_r<33> a_blc_r<32> a_blt_r<35> a_blt_r<34> a_blt_r<33> a_blt_r<32> A_BM<40> a_dclk_n_r<8> a_dclk_n_r<9> a_dclk_p_r<8> a_dclk_p_r<9> A_DOUT<40> A_DIN<40> a_rclk_n_r<8> a_rclk_n_r<9> a_rclk_p_r<8> a_rclk_p_r<9> a_tieh<40> a_wclk_n_r<8> a_wclk_n_r<9> a_wclk_p_r<8> a_wclk_p_r<9> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<39> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<39> A_BIST_DIN<39> A_BIST_EN a_blc_r<31> a_blc_r<30> a_blc_r<29> a_blc_r<28> a_blt_r<31> a_blt_r<30> a_blt_r<29> a_blt_r<28> A_BM<39> a_dclk_n_r<7> a_dclk_n_r<8> a_dclk_p_r<7> a_dclk_p_r<8> A_DOUT<39> A_DIN<39> a_rclk_n_r<7> a_rclk_n_r<8> a_rclk_p_r<7> a_rclk_p_r<8> a_tieh<39> a_wclk_n_r<7> a_wclk_n_r<8> a_wclk_p_r<7> a_wclk_p_r<8> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<38> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<38> A_BIST_DIN<38> A_BIST_EN a_blc_r<27> a_blc_r<26> a_blc_r<25> a_blc_r<24> a_blt_r<27> a_blt_r<26> a_blt_r<25> a_blt_r<24> A_BM<38> a_dclk_n_r<6> a_dclk_n_r<7> a_dclk_p_r<6> a_dclk_p_r<7> A_DOUT<38> A_DIN<38> a_rclk_n_r<6> a_rclk_n_r<7> a_rclk_p_r<6> a_rclk_p_r<7> a_tieh<38> a_wclk_n_r<6> a_wclk_n_r<7> a_wclk_p_r<6> a_wclk_p_r<7> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<37> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<37> A_BIST_DIN<37> A_BIST_EN a_blc_r<23> a_blc_r<22> a_blc_r<21> a_blc_r<20> a_blt_r<23> a_blt_r<22> a_blt_r<21> a_blt_r<20> A_BM<37> a_dclk_n_r<5> a_dclk_n_r<6> a_dclk_p_r<5> a_dclk_p_r<6> A_DOUT<37> A_DIN<37> a_rclk_n_r<5> a_rclk_n_r<6> a_rclk_p_r<5> a_rclk_p_r<6> a_tieh<37> a_wclk_n_r<5> a_wclk_n_r<6> a_wclk_p_r<5> a_wclk_p_r<6> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<36> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<36> A_BIST_DIN<36> A_BIST_EN a_blc_r<19> a_blc_r<18> a_blc_r<17> a_blc_r<16> a_blt_r<19> a_blt_r<18> a_blt_r<17> a_blt_r<16> A_BM<36> a_dclk_n_r<4> a_dclk_n_r<5> a_dclk_p_r<4> a_dclk_p_r<5> A_DOUT<36> A_DIN<36> a_rclk_n_r<4> a_rclk_n_r<5> a_rclk_p_r<4> a_rclk_p_r<5> a_tieh<36> a_wclk_n_r<4> a_wclk_n_r<5> a_wclk_p_r<4> a_wclk_p_r<5> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<35> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<35> A_BIST_DIN<35> A_BIST_EN a_blc_r<15> a_blc_r<14> a_blc_r<13> a_blc_r<12> a_blt_r<15> a_blt_r<14> a_blt_r<13> a_blt_r<12> A_BM<35> a_dclk_n_r<3> a_dclk_n_r<4> a_dclk_p_r<3> a_dclk_p_r<4> A_DOUT<35> A_DIN<35> a_rclk_n_r<3> a_rclk_n_r<4> a_rclk_p_r<3> a_rclk_p_r<4> a_tieh<35> a_wclk_n_r<3> a_wclk_n_r<4> a_wclk_p_r<3> a_wclk_p_r<4> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<34> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<34> A_BIST_DIN<34> A_BIST_EN a_blc_r<11> a_blc_r<10> a_blc_r<9> a_blc_r<8> a_blt_r<11> a_blt_r<10> a_blt_r<9> a_blt_r<8> A_BM<34> a_dclk_n_r<2> a_dclk_n_r<3> a_dclk_p_r<2> a_dclk_p_r<3> A_DOUT<34> A_DIN<34> a_rclk_n_r<2> a_rclk_n_r<3> a_rclk_p_r<2> a_rclk_p_r<3> a_tieh<34> a_wclk_n_r<2> a_wclk_n_r<3> a_wclk_p_r<2> a_wclk_p_r<3> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<33> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<33> A_BIST_DIN<33> A_BIST_EN a_blc_r<7> a_blc_r<6> a_blc_r<5> a_blc_r<4> a_blt_r<7> a_blt_r<6> a_blt_r<5> a_blt_r<4> A_BM<33> a_dclk_n_r<1> a_dclk_n_r<2> a_dclk_p_r<1> a_dclk_p_r<2> A_DOUT<33> A_DIN<33> a_rclk_n_r<1> a_rclk_n_r<2> a_rclk_p_r<1> a_rclk_p_r<2> a_tieh<33> a_wclk_n_r<1> a_wclk_n_r<2> a_wclk_p_r<1> a_wclk_p_r<2> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<32> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<32> A_BIST_DIN<32> A_BIST_EN a_blc_r<3> a_blc_r<2> a_blc_r<1> a_blc_r<0> a_blt_r<3> a_blt_r<2> a_blt_r<1> a_blt_r<0> A_BM<32> a_dclk_n_r<0> a_dclk_n_r<1> a_dclk_p_r<0> a_dclk_p_r<1> A_DOUT<32> A_DIN<32> a_rclk_n_r<0> a_rclk_n_r<1> a_rclk_p_r<0> a_rclk_p_r<1> a_tieh<32> a_wclk_n_r<0> a_wclk_n_r<1> a_wclk_p_r<0> a_wclk_p_r<1> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<31> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<0> A_BIST_DIN<0> A_BIST_EN a_blc_l<127> a_blc_l<126> a_blc_l<125> a_blc_l<124> a_blt_l<127> a_blt_l<126> a_blt_l<125> a_blt_l<124> A_BM<0> a_dclk_n_l<31> a_dclk_n_l<32> a_dclk_p_l<31> a_dclk_p_l<32> A_DOUT<0> A_DIN<0> a_rclk_n_l<31> a_rclk_n_l<32> a_rclk_p_l<31> a_rclk_p_l<32> a_tieh<0> a_wclk_n_l<31> a_wclk_n_l<32> a_wclk_p_l<31> a_wclk_p_l<32> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<30> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<1> A_BIST_DIN<1> A_BIST_EN a_blc_l<123> a_blc_l<122> a_blc_l<121> a_blc_l<120> a_blt_l<123> a_blt_l<122> a_blt_l<121> a_blt_l<120> A_BM<1> a_dclk_n_l<30> a_dclk_n_l<31> a_dclk_p_l<30> a_dclk_p_l<31> A_DOUT<1> A_DIN<1> a_rclk_n_l<30> a_rclk_n_l<31> a_rclk_p_l<30> a_rclk_p_l<31> a_tieh<1> a_wclk_n_l<30> a_wclk_n_l<31> a_wclk_p_l<30> a_wclk_p_l<31> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<29> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<2> A_BIST_DIN<2> A_BIST_EN a_blc_l<119> a_blc_l<118> a_blc_l<117> a_blc_l<116> a_blt_l<119> a_blt_l<118> a_blt_l<117> a_blt_l<116> A_BM<2> a_dclk_n_l<29> a_dclk_n_l<30> a_dclk_p_l<29> a_dclk_p_l<30> A_DOUT<2> A_DIN<2> a_rclk_n_l<29> a_rclk_n_l<30> a_rclk_p_l<29> a_rclk_p_l<30> a_tieh<2> a_wclk_n_l<29> a_wclk_n_l<30> a_wclk_p_l<29> a_wclk_p_l<30> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<28> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<3> A_BIST_DIN<3> A_BIST_EN a_blc_l<115> a_blc_l<114> a_blc_l<113> a_blc_l<112> a_blt_l<115> a_blt_l<114> a_blt_l<113> a_blt_l<112> A_BM<3> a_dclk_n_l<28> a_dclk_n_l<29> a_dclk_p_l<28> a_dclk_p_l<29> A_DOUT<3> A_DIN<3> a_rclk_n_l<28> a_rclk_n_l<29> a_rclk_p_l<28> a_rclk_p_l<29> a_tieh<3> a_wclk_n_l<28> a_wclk_n_l<29> a_wclk_p_l<28> a_wclk_p_l<29> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<27> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<4> A_BIST_DIN<4> A_BIST_EN a_blc_l<111> a_blc_l<110> a_blc_l<109> a_blc_l<108> a_blt_l<111> a_blt_l<110> a_blt_l<109> a_blt_l<108> A_BM<4> a_dclk_n_l<27> a_dclk_n_l<28> a_dclk_p_l<27> a_dclk_p_l<28> A_DOUT<4> A_DIN<4> a_rclk_n_l<27> a_rclk_n_l<28> a_rclk_p_l<27> a_rclk_p_l<28> a_tieh<4> a_wclk_n_l<27> a_wclk_n_l<28> a_wclk_p_l<27> a_wclk_p_l<28> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<26> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<5> A_BIST_DIN<5> A_BIST_EN a_blc_l<107> a_blc_l<106> a_blc_l<105> a_blc_l<104> a_blt_l<107> a_blt_l<106> a_blt_l<105> a_blt_l<104> A_BM<5> a_dclk_n_l<26> a_dclk_n_l<27> a_dclk_p_l<26> a_dclk_p_l<27> A_DOUT<5> A_DIN<5> a_rclk_n_l<26> a_rclk_n_l<27> a_rclk_p_l<26> a_rclk_p_l<27> a_tieh<5> a_wclk_n_l<26> a_wclk_n_l<27> a_wclk_p_l<26> a_wclk_p_l<27> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<25> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<6> A_BIST_DIN<6> A_BIST_EN a_blc_l<103> a_blc_l<102> a_blc_l<101> a_blc_l<100> a_blt_l<103> a_blt_l<102> a_blt_l<101> a_blt_l<100> A_BM<6> a_dclk_n_l<25> a_dclk_n_l<26> a_dclk_p_l<25> a_dclk_p_l<26> A_DOUT<6> A_DIN<6> a_rclk_n_l<25> a_rclk_n_l<26> a_rclk_p_l<25> a_rclk_p_l<26> a_tieh<6> a_wclk_n_l<25> a_wclk_n_l<26> a_wclk_p_l<25> a_wclk_p_l<26> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<24> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<7> A_BIST_DIN<7> A_BIST_EN a_blc_l<99> a_blc_l<98> a_blc_l<97> a_blc_l<96> a_blt_l<99> a_blt_l<98> a_blt_l<97> a_blt_l<96> A_BM<7> a_dclk_n_l<24> a_dclk_n_l<25> a_dclk_p_l<24> a_dclk_p_l<25> A_DOUT<7> A_DIN<7> a_rclk_n_l<24> a_rclk_n_l<25> a_rclk_p_l<24> a_rclk_p_l<25> a_tieh<7> a_wclk_n_l<24> a_wclk_n_l<25> a_wclk_p_l<24> a_wclk_p_l<25> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<23> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<8> A_BIST_DIN<8> A_BIST_EN a_blc_l<95> a_blc_l<94> a_blc_l<93> a_blc_l<92> a_blt_l<95> a_blt_l<94> a_blt_l<93> a_blt_l<92> A_BM<8> a_dclk_n_l<23> a_dclk_n_l<24> a_dclk_p_l<23> a_dclk_p_l<24> A_DOUT<8> A_DIN<8> a_rclk_n_l<23> a_rclk_n_l<24> a_rclk_p_l<23> a_rclk_p_l<24> a_tieh<8> a_wclk_n_l<23> a_wclk_n_l<24> a_wclk_p_l<23> a_wclk_p_l<24> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<22> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<9> A_BIST_DIN<9> A_BIST_EN a_blc_l<91> a_blc_l<90> a_blc_l<89> a_blc_l<88> a_blt_l<91> a_blt_l<90> a_blt_l<89> a_blt_l<88> A_BM<9> a_dclk_n_l<22> a_dclk_n_l<23> a_dclk_p_l<22> a_dclk_p_l<23> A_DOUT<9> A_DIN<9> a_rclk_n_l<22> a_rclk_n_l<23> a_rclk_p_l<22> a_rclk_p_l<23> a_tieh<9> a_wclk_n_l<22> a_wclk_n_l<23> a_wclk_p_l<22> a_wclk_p_l<23> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<21> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<10> A_BIST_DIN<10> A_BIST_EN a_blc_l<87> a_blc_l<86> a_blc_l<85> a_blc_l<84> a_blt_l<87> a_blt_l<86> a_blt_l<85> a_blt_l<84> A_BM<10> a_dclk_n_l<21> a_dclk_n_l<22> a_dclk_p_l<21> a_dclk_p_l<22> A_DOUT<10> A_DIN<10> a_rclk_n_l<21> a_rclk_n_l<22> a_rclk_p_l<21> a_rclk_p_l<22> a_tieh<10> a_wclk_n_l<21> a_wclk_n_l<22> a_wclk_p_l<21> a_wclk_p_l<22> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<20> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<11> A_BIST_DIN<11> A_BIST_EN a_blc_l<83> a_blc_l<82> a_blc_l<81> a_blc_l<80> a_blt_l<83> a_blt_l<82> a_blt_l<81> a_blt_l<80> A_BM<11> a_dclk_n_l<20> a_dclk_n_l<21> a_dclk_p_l<20> a_dclk_p_l<21> A_DOUT<11> A_DIN<11> a_rclk_n_l<20> a_rclk_n_l<21> a_rclk_p_l<20> a_rclk_p_l<21> a_tieh<11> a_wclk_n_l<20> a_wclk_n_l<21> a_wclk_p_l<20> a_wclk_p_l<21> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<19> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<12> A_BIST_DIN<12> A_BIST_EN a_blc_l<79> a_blc_l<78> a_blc_l<77> a_blc_l<76> a_blt_l<79> a_blt_l<78> a_blt_l<77> a_blt_l<76> A_BM<12> a_dclk_n_l<19> a_dclk_n_l<20> a_dclk_p_l<19> a_dclk_p_l<20> A_DOUT<12> A_DIN<12> a_rclk_n_l<19> a_rclk_n_l<20> a_rclk_p_l<19> a_rclk_p_l<20> a_tieh<12> a_wclk_n_l<19> a_wclk_n_l<20> a_wclk_p_l<19> a_wclk_p_l<20> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<18> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<13> A_BIST_DIN<13> A_BIST_EN a_blc_l<75> a_blc_l<74> a_blc_l<73> a_blc_l<72> a_blt_l<75> a_blt_l<74> a_blt_l<73> a_blt_l<72> A_BM<13> a_dclk_n_l<18> a_dclk_n_l<19> a_dclk_p_l<18> a_dclk_p_l<19> A_DOUT<13> A_DIN<13> a_rclk_n_l<18> a_rclk_n_l<19> a_rclk_p_l<18> a_rclk_p_l<19> a_tieh<13> a_wclk_n_l<18> a_wclk_n_l<19> a_wclk_p_l<18> a_wclk_p_l<19> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<17> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<14> A_BIST_DIN<14> A_BIST_EN a_blc_l<71> a_blc_l<70> a_blc_l<69> a_blc_l<68> a_blt_l<71> a_blt_l<70> a_blt_l<69> a_blt_l<68> A_BM<14> a_dclk_n_l<17> a_dclk_n_l<18> a_dclk_p_l<17> a_dclk_p_l<18> A_DOUT<14> A_DIN<14> a_rclk_n_l<17> a_rclk_n_l<18> a_rclk_p_l<17> a_rclk_p_l<18> a_tieh<14> a_wclk_n_l<17> a_wclk_n_l<18> a_wclk_p_l<17> a_wclk_p_l<18> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<16> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<15> A_BIST_DIN<15> A_BIST_EN a_blc_l<67> a_blc_l<66> a_blc_l<65> a_blc_l<64> a_blt_l<67> a_blt_l<66> a_blt_l<65> a_blt_l<64> A_BM<15> a_dclk_n_l<16> a_dclk_n_l<17> a_dclk_p_l<16> a_dclk_p_l<17> A_DOUT<15> A_DIN<15> a_rclk_n_l<16> a_rclk_n_l<17> a_rclk_p_l<16> a_rclk_p_l<17> a_tieh<15> a_wclk_n_l<16> a_wclk_n_l<17> a_wclk_p_l<16> a_wclk_p_l<17> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<15> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<16> A_BIST_DIN<16> A_BIST_EN a_blc_l<63> a_blc_l<62> a_blc_l<61> a_blc_l<60> a_blt_l<63> a_blt_l<62> a_blt_l<61> a_blt_l<60> A_BM<16> a_dclk_n_l<15> a_dclk_n_l<16> a_dclk_p_l<15> a_dclk_p_l<16> A_DOUT<16> A_DIN<16> a_rclk_n_l<15> a_rclk_n_l<16> a_rclk_p_l<15> a_rclk_p_l<16> a_tieh<16> a_wclk_n_l<15> a_wclk_n_l<16> a_wclk_p_l<15> a_wclk_p_l<16> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<14> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<17> A_BIST_DIN<17> A_BIST_EN a_blc_l<59> a_blc_l<58> a_blc_l<57> a_blc_l<56> a_blt_l<59> a_blt_l<58> a_blt_l<57> a_blt_l<56> A_BM<17> a_dclk_n_l<14> a_dclk_n_l<15> a_dclk_p_l<14> a_dclk_p_l<15> A_DOUT<17> A_DIN<17> a_rclk_n_l<14> a_rclk_n_l<15> a_rclk_p_l<14> a_rclk_p_l<15> a_tieh<17> a_wclk_n_l<14> a_wclk_n_l<15> a_wclk_p_l<14> a_wclk_p_l<15> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<13> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<18> A_BIST_DIN<18> A_BIST_EN a_blc_l<55> a_blc_l<54> a_blc_l<53> a_blc_l<52> a_blt_l<55> a_blt_l<54> a_blt_l<53> a_blt_l<52> A_BM<18> a_dclk_n_l<13> a_dclk_n_l<14> a_dclk_p_l<13> a_dclk_p_l<14> A_DOUT<18> A_DIN<18> a_rclk_n_l<13> a_rclk_n_l<14> a_rclk_p_l<13> a_rclk_p_l<14> a_tieh<18> a_wclk_n_l<13> a_wclk_n_l<14> a_wclk_p_l<13> a_wclk_p_l<14> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<12> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<19> A_BIST_DIN<19> A_BIST_EN a_blc_l<51> a_blc_l<50> a_blc_l<49> a_blc_l<48> a_blt_l<51> a_blt_l<50> a_blt_l<49> a_blt_l<48> A_BM<19> a_dclk_n_l<12> a_dclk_n_l<13> a_dclk_p_l<12> a_dclk_p_l<13> A_DOUT<19> A_DIN<19> a_rclk_n_l<12> a_rclk_n_l<13> a_rclk_p_l<12> a_rclk_p_l<13> a_tieh<19> a_wclk_n_l<12> a_wclk_n_l<13> a_wclk_p_l<12> a_wclk_p_l<13> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<11> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<20> A_BIST_DIN<20> A_BIST_EN a_blc_l<47> a_blc_l<46> a_blc_l<45> a_blc_l<44> a_blt_l<47> a_blt_l<46> a_blt_l<45> a_blt_l<44> A_BM<20> a_dclk_n_l<11> a_dclk_n_l<12> a_dclk_p_l<11> a_dclk_p_l<12> A_DOUT<20> A_DIN<20> a_rclk_n_l<11> a_rclk_n_l<12> a_rclk_p_l<11> a_rclk_p_l<12> a_tieh<20> a_wclk_n_l<11> a_wclk_n_l<12> a_wclk_p_l<11> a_wclk_p_l<12> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<10> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<21> A_BIST_DIN<21> A_BIST_EN a_blc_l<43> a_blc_l<42> a_blc_l<41> a_blc_l<40> a_blt_l<43> a_blt_l<42> a_blt_l<41> a_blt_l<40> A_BM<21> a_dclk_n_l<10> a_dclk_n_l<11> a_dclk_p_l<10> a_dclk_p_l<11> A_DOUT<21> A_DIN<21> a_rclk_n_l<10> a_rclk_n_l<11> a_rclk_p_l<10> a_rclk_p_l<11> a_tieh<21> a_wclk_n_l<10> a_wclk_n_l<11> a_wclk_p_l<10> a_wclk_p_l<11> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<9> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<22> A_BIST_DIN<22> A_BIST_EN a_blc_l<39> a_blc_l<38> a_blc_l<37> a_blc_l<36> a_blt_l<39> a_blt_l<38> a_blt_l<37> a_blt_l<36> A_BM<22> a_dclk_n_l<9> a_dclk_n_l<10> a_dclk_p_l<9> a_dclk_p_l<10> A_DOUT<22> A_DIN<22> a_rclk_n_l<9> a_rclk_n_l<10> a_rclk_p_l<9> a_rclk_p_l<10> a_tieh<22> a_wclk_n_l<9> a_wclk_n_l<10> a_wclk_p_l<9> a_wclk_p_l<10> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<8> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<23> A_BIST_DIN<23> A_BIST_EN a_blc_l<35> a_blc_l<34> a_blc_l<33> a_blc_l<32> a_blt_l<35> a_blt_l<34> a_blt_l<33> a_blt_l<32> A_BM<23> a_dclk_n_l<8> a_dclk_n_l<9> a_dclk_p_l<8> a_dclk_p_l<9> A_DOUT<23> A_DIN<23> a_rclk_n_l<8> a_rclk_n_l<9> a_rclk_p_l<8> a_rclk_p_l<9> a_tieh<23> a_wclk_n_l<8> a_wclk_n_l<9> a_wclk_p_l<8> a_wclk_p_l<9> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<7> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<24> A_BIST_DIN<24> A_BIST_EN a_blc_l<31> a_blc_l<30> a_blc_l<29> a_blc_l<28> a_blt_l<31> a_blt_l<30> a_blt_l<29> a_blt_l<28> A_BM<24> a_dclk_n_l<7> a_dclk_n_l<8> a_dclk_p_l<7> a_dclk_p_l<8> A_DOUT<24> A_DIN<24> a_rclk_n_l<7> a_rclk_n_l<8> a_rclk_p_l<7> a_rclk_p_l<8> a_tieh<24> a_wclk_n_l<7> a_wclk_n_l<8> a_wclk_p_l<7> a_wclk_p_l<8> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<6> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<25> A_BIST_DIN<25> A_BIST_EN a_blc_l<27> a_blc_l<26> a_blc_l<25> a_blc_l<24> a_blt_l<27> a_blt_l<26> a_blt_l<25> a_blt_l<24> A_BM<25> a_dclk_n_l<6> a_dclk_n_l<7> a_dclk_p_l<6> a_dclk_p_l<7> A_DOUT<25> A_DIN<25> a_rclk_n_l<6> a_rclk_n_l<7> a_rclk_p_l<6> a_rclk_p_l<7> a_tieh<25> a_wclk_n_l<6> a_wclk_n_l<7> a_wclk_p_l<6> a_wclk_p_l<7> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<5> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<26> A_BIST_DIN<26> A_BIST_EN a_blc_l<23> a_blc_l<22> a_blc_l<21> a_blc_l<20> a_blt_l<23> a_blt_l<22> a_blt_l<21> a_blt_l<20> A_BM<26> a_dclk_n_l<5> a_dclk_n_l<6> a_dclk_p_l<5> a_dclk_p_l<6> A_DOUT<26> A_DIN<26> a_rclk_n_l<5> a_rclk_n_l<6> a_rclk_p_l<5> a_rclk_p_l<6> a_tieh<26> a_wclk_n_l<5> a_wclk_n_l<6> a_wclk_p_l<5> a_wclk_p_l<6> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<4> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<27> A_BIST_DIN<27> A_BIST_EN a_blc_l<19> a_blc_l<18> a_blc_l<17> a_blc_l<16> a_blt_l<19> a_blt_l<18> a_blt_l<17> a_blt_l<16> A_BM<27> a_dclk_n_l<4> a_dclk_n_l<5> a_dclk_p_l<4> a_dclk_p_l<5> A_DOUT<27> A_DIN<27> a_rclk_n_l<4> a_rclk_n_l<5> a_rclk_p_l<4> a_rclk_p_l<5> a_tieh<27> a_wclk_n_l<4> a_wclk_n_l<5> a_wclk_p_l<4> a_wclk_p_l<5> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<3> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<28> A_BIST_DIN<28> A_BIST_EN a_blc_l<15> a_blc_l<14> a_blc_l<13> a_blc_l<12> a_blt_l<15> a_blt_l<14> a_blt_l<13> a_blt_l<12> A_BM<28> a_dclk_n_l<3> a_dclk_n_l<4> a_dclk_p_l<3> a_dclk_p_l<4> A_DOUT<28> A_DIN<28> a_rclk_n_l<3> a_rclk_n_l<4> a_rclk_p_l<3> a_rclk_p_l<4> a_tieh<28> a_wclk_n_l<3> a_wclk_n_l<4> a_wclk_p_l<3> a_wclk_p_l<4> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<2> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<29> A_BIST_DIN<29> A_BIST_EN a_blc_l<11> a_blc_l<10> a_blc_l<9> a_blc_l<8> a_blt_l<11> a_blt_l<10> a_blt_l<9> a_blt_l<8> A_BM<29> a_dclk_n_l<2> a_dclk_n_l<3> a_dclk_p_l<2> a_dclk_p_l<3> A_DOUT<29> A_DIN<29> a_rclk_n_l<2> a_rclk_n_l<3> a_rclk_p_l<2> a_rclk_p_l<3> a_tieh<29> a_wclk_n_l<2> a_wclk_n_l<3> a_wclk_p_l<2> a_wclk_p_l<3> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<1> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<30> A_BIST_DIN<30> A_BIST_EN a_blc_l<7> a_blc_l<6> a_blc_l<5> a_blc_l<4> a_blt_l<7> a_blt_l<6> a_blt_l<5> a_blt_l<4> A_BM<30> a_dclk_n_l<1> a_dclk_n_l<2> a_dclk_p_l<1> a_dclk_p_l<2> A_DOUT<30> A_DIN<30> a_rclk_n_l<1> a_rclk_n_l<2> a_rclk_p_l<1> a_rclk_p_l<2> a_tieh<30> a_wclk_n_l<1> a_wclk_n_l<2> a_wclk_p_l<1> a_wclk_p_l<2> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2
XCOLCTRL<0> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<31> A_BIST_DIN<31> A_BIST_EN a_blc_l<3> a_blc_l<2> a_blc_l<1> a_blc_l<0> a_blt_l<3> a_blt_l<2> a_blt_l<1> a_blt_l<0> A_BM<31> a_dclk_n_l<0> a_dclk_n_l<1> a_dclk_p_l<0> a_dclk_p_l<1> A_DOUT<31> A_DIN<31> a_rclk_n_l<0> a_rclk_n_l<1> a_rclk_p_l<0> a_rclk_p_l<1> a_tieh<31> a_wclk_n_l<0> a_wclk_n_l<1> a_wclk_p_l<0> a_wclk_p_l<1> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLCTRL2


XDRVFILL4<1> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4
XDRVFILL4<2> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4
XDRVFILL4<3> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4
XDRVFILL4<4> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4
XCOLFILL4<1> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<2> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<3> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<4> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<5> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<6> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<7> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<8> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<9> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<10> VDD! VSS! / RM_IHPSG13_1024x64_c2_1P_COLDRV13_FILL4C2
.ENDS
