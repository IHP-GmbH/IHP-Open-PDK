************************************************************************
* 
* Copyright 2023 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
************************************************************************

.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_CORNER VDD_CORE VSS
XI16 VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR LWL NW PW VDD VSS
MN1 VSS LWL VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 VSS net9 VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR A_WL<15> A_WL<14> A_WL<13> A_WL<12> 
+ A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> 
+ A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS
XI0<15> A_WL<15> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<14> A_WL<14> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<13> A_WL<13> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<12> A_WL<12> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<11> A_WL<11> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<10> A_WL<10> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<9> A_WL<9> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<8> A_WL<8> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<7> A_WL<7> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<6> A_WL<6> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<5> A_WL<5> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<4> A_WL<4> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<3> A_WL<3> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<2> A_WL<2> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<1> A_WL<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
XI0<0> A_WL<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_LR
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL BLC_BOT BLC_TOP BLT_BOT BLT_TOP LWL NW PW 
+ RWL VDD VSS
MN0 NC NT VSS PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN1 NT NC VSS PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN3 NC RWL BLC_TOP PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN2 BLT_BOT LWL NT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 NT NC VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 NC NT VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
R1 BLC_BOT BLC_TOP lvsres w=2.6e-07 l=6e-07
R0 BLT_BOT BLT_TOP lvsres w=2.6e-07 l=6e-07
R2 RWL LWL lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> 
+ A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<15> 
+ A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> 
+ A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> 
+ A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> 
+ A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE 
+ VSS
XCELL<31> A_BLC_TOP<1> A_RBLC<15> A_BLT_TOP<1> A_RBLT<15> A_RWL<15> 
+ VDD_CORE VSS A_XWL<15> VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<30> A_RBLC<14> A_RBLC<15> A_RBLT<14> A_RBLT<15> A_RWL<14> VDD_CORE 
+ VSS A_XWL<14> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<29> A_RBLC<14> A_RBLC<13> A_RBLT<14> A_RBLT<13> A_RWL<13> VDD_CORE 
+ VSS A_XWL<13> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<28> A_RBLC<12> A_RBLC<13> A_RBLT<12> A_RBLT<13> A_RWL<12> VDD_CORE 
+ VSS A_XWL<12> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<27> A_RBLC<12> A_RBLC<11> A_RBLT<12> A_RBLT<11> A_RWL<11> VDD_CORE 
+ VSS A_XWL<11> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<26> A_RBLC<10> A_RBLC<11> A_RBLT<10> A_RBLT<11> A_RWL<10> VDD_CORE 
+ VSS A_XWL<10> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<25> A_RBLC<10> A_RBLC<9> A_RBLT<10> A_RBLT<9> A_RWL<9> VDD_CORE 
+ VSS A_XWL<9> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<24> A_RBLC<8> A_RBLC<9> A_RBLT<8> A_RBLT<9> A_RWL<8> VDD_CORE 
+ VSS A_XWL<8> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<23> A_RBLC<8> A_RBLC<7> A_RBLT<8> A_RBLT<7> A_RWL<7> VDD_CORE 
+ VSS A_XWL<7> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<22> A_RBLC<6> A_RBLC<7> A_RBLT<6> A_RBLT<7> A_RWL<6> VDD_CORE 
+ VSS A_XWL<6> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<21> A_RBLC<6> A_RBLC<5> A_RBLT<6> A_RBLT<5> A_RWL<5> VDD_CORE 
+ VSS A_XWL<5> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<20> A_RBLC<4> A_RBLC<5> A_RBLT<4> A_RBLT<5> A_RWL<4> VDD_CORE 
+ VSS A_XWL<4> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<19> A_RBLC<4> A_RBLC<3> A_RBLT<4> A_RBLT<3> A_RWL<3> VDD_CORE 
+ VSS A_XWL<3> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<18> A_RBLC<2> A_RBLC<3> A_RBLT<2> A_RBLT<3> A_RWL<2> VDD_CORE 
+ VSS A_XWL<2> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<17> A_RBLC<2> A_RBLC<1> A_RBLT<2> A_RBLT<1> A_RWL<1> VDD_CORE 
+ VSS A_XWL<1> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<16> A_BLC_BOT<1> A_RBLC<1> A_BLT_BOT<1> A_RBLT<1> A_RWL<0> VDD_CORE 
+ VSS A_XWL<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<15> A_BLC_TOP<0> A_LBLC<15> A_BLT_TOP<0> A_LBLT<15> A_LWL<15> 
+ VDD_CORE VSS A_XWL<15> VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<14> A_LBLC<14> A_LBLC<15> A_LBLT<14> A_LBLT<15> A_LWL<14> VDD_CORE 
+ VSS A_XWL<14> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<13> A_LBLC<14> A_LBLC<13> A_LBLT<14> A_LBLT<13> A_LWL<13> VDD_CORE 
+ VSS A_XWL<13> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<12> A_LBLC<12> A_LBLC<13> A_LBLT<12> A_LBLT<13> A_LWL<12> VDD_CORE 
+ VSS A_XWL<12> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<11> A_LBLC<12> A_LBLC<11> A_LBLT<12> A_LBLT<11> A_LWL<11> VDD_CORE 
+ VSS A_XWL<11> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<10> A_LBLC<10> A_LBLC<11> A_LBLT<10> A_LBLT<11> A_LWL<10> VDD_CORE 
+ VSS A_XWL<10> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<9> A_LBLC<10> A_LBLC<9> A_LBLT<10> A_LBLT<9> A_LWL<9> VDD_CORE 
+ VSS A_XWL<9> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<8> A_LBLC<8> A_LBLC<9> A_LBLT<8> A_LBLT<9> A_LWL<8> VDD_CORE 
+ VSS A_XWL<8> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<7> A_LBLC<8> A_LBLC<7> A_LBLT<8> A_LBLT<7> A_LWL<7> VDD_CORE 
+ VSS A_XWL<7> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<6> A_LBLC<6> A_LBLC<7> A_LBLT<6> A_LBLT<7> A_LWL<6> VDD_CORE 
+ VSS A_XWL<6> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<5> A_LBLC<6> A_LBLC<5> A_LBLT<6> A_LBLT<5> A_LWL<5> VDD_CORE 
+ VSS A_XWL<5> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<4> A_LBLC<4> A_LBLC<5> A_LBLT<4> A_LBLT<5> A_LWL<4> VDD_CORE 
+ VSS A_XWL<4> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<3> A_LBLC<4> A_LBLC<3> A_LBLT<4> A_LBLT<3> A_LWL<3> VDD_CORE 
+ VSS A_XWL<3> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<2> A_LBLC<2> A_LBLC<3> A_LBLT<2> A_LBLT<3> A_LWL<2> VDD_CORE 
+ VSS A_XWL<2> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<1> A_LBLC<2> A_LBLC<1> A_LBLT<2> A_LBLT<1> A_LWL<1> VDD_CORE 
+ VSS A_XWL<1> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
XCELL<0> A_BLC_BOT<0> A_LBLC<1> A_BLT_BOT<0> A_LBLT<1> A_LWL<0> VDD_CORE 
+ VSS A_XWL<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_CELL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB BLC BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_TB A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ VDD_CORE VSS
XEDGE<1> A_BLC<1> A_BLT<1> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB
XEDGE<0> A_BLC<0> A_BLT<0> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB
.ENDS

.SUBCKT RSC_IHPSG13_CBUFX4 A Z VDD VSS
MN0 net9 A VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 Z net9 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP0 net9 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 Z net9 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDRV13X4 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX4 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net6 A VSS VSS nmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_WLDRV16X4 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX4
.ENDS
.SUBCKT RSC_IHPSG13_FILLCAP8 VDD VSS
MN0 vss_r vdd_r VSS VSS nmos m=1 w=4.98u l=130.00n ng=6 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD pmos m=1 w=6.48u l=385.000n ng=4 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_LHPQX2 CP D Q VDD VSS
MN3 QIN CPN net14 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN2 net14 net10 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN5 net21 D VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 QIN CP net21 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net10 QIN VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 CPN CP VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 Q QIN VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP2 QIN CP net16 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 CPN CP VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 Q QIN VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP3 net10 QIN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net16 net10 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP6 QIN CPN net20 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP5 net20 D VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NAND2X2 A B Z VDD VSS
MP1 Z B VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN0 Z B net7 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net7 A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX4 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX2 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_INVX2 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NAND3X2 A B C Z VDD VSS
MP2 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 Z B VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z C VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN1 net12 B net16 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN0 Z C net12 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN2 net16 A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_NOR3X2 A B C Z VDD VSS
MP0 net13 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP2 Z C net10 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP1 net10 B net13 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN1 Z B VSS VSS nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
MN0 Z C VSS VSS nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
MN2 Z A VSS VSS nmos m=1 w=875.000n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_FILLCAP4 VDD VSS
MN0 vss_r vdd_r VSS VSS nmos m=1 w=2.49u l=130.00n ng=3 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD pmos m=1 w=3.24u l=385.000n ng=2 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MET2RES A B
R0 B A lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_DEC04 ADDR<3> ADDR<2> ADDR<1> ADDR<0> CS ECLK_H_BOT 
+ ECLK_H_TOP ECLK_L_BOT ECLK_L_TOP WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> 
+ WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> VDD VSS
XLATCH<3> CS ADDR<3> PADR<3> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<2> CS ADDR<2> PADR<2> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<1> CS ADDR<1> PADR<1> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<0> CS ADDR<0> PADR<0> VDD VSS / RSC_IHPSG13_LHPQX2
XI0<3> PADR<1> PADR<0> sel01<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<2> PADR<1> NADR<0> sel01<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<1> NADR<1> PADR<0> sel01<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<0> NADR<1> NADR<0> sel01<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI4 ECLK_L_BOT EN VDD VSS / RSC_IHPSG13_CINVX4
XI5 ECLK_H_BOT ECLK_L_BOT VDD VSS / RSC_IHPSG13_CINVX2
XI3<3> PADR<3> NADR<3> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> PADR<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> PADR<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> PADR<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1<3> PADR<2> PADR<3> CS sel23<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<2> PADR<3> CS sel23<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<2> NADR<3> CS sel23<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<2> NADR<3> CS sel23<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI2<15> sel23<3> sel01<3> EN WL<15> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<14> sel23<3> sel01<2> EN WL<14> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<13> sel23<3> sel01<1> EN WL<13> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<12> sel23<3> sel01<0> EN WL<12> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<11> sel23<2> sel01<3> EN WL<11> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<10> sel23<2> sel01<2> EN WL<10> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<9> sel23<2> sel01<1> EN WL<9> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<8> sel23<2> sel01<0> EN WL<8> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<7> sel23<1> sel01<3> EN WL<7> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<6> sel23<1> sel01<2> EN WL<6> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<5> sel23<1> sel01<1> EN WL<5> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<4> sel23<1> sel01<0> EN WL<4> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<3> sel23<0> sel01<3> EN WL<3> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<2> sel23<0> sel01<2> EN WL<2> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<1> sel23<0> sel01<1> EN WL<1> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<0> sel23<0> sel01<0> EN WL<0> VDD VSS / RSC_IHPSG13_NOR3X2
XCAPS4 VDD VSS / RSC_IHPSG13_FILLCAP4
XI11 ECLK_L_BOT ECLK_L_TOP / RSC_IHPSG13_MET2RES
XR0 ECLK_H_BOT ECLK_H_TOP / RSC_IHPSG13_MET2RES
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWDEC4 ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> 
+ CS_I ECLK_I WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XSEL ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I ECLK_H<1> 
+ ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> 
+ WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> 
+ WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
.ENDS
.SUBCKT RSC_IHPSG13_CINVX8 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=2.82u l=130.00n ng=4 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_DFNQMX2IX1 BE BI CN D QI QIN VDD VSS
MN15 net026 BI VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN14 MXI_OUT BE net026 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net025 D VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 MXI_OUT BEN net025 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN10 QI CNN net21 VSS nmos m=1 w=850.00n l=130.00n ng=1 nrd=0 nrs=0
MN11 net21 QI_MS VSS VSS nmos m=1 w=850.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN7 net30 QI_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN6 QIN_MS CNN net30 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 QI_MS QIN_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN12 CNN CN VSS VSS nmos m=1 w=495.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN9 net37 MXI_OUT VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN8 QIN_MS CN net37 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 QI CN net25 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN4 net25 QIN VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 QIN QI VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN13 BEN BE VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP15 MXI_OUT BEN net027 VDD pmos m=1 w=985.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP14 net027 BI VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP1 MXI_OUT BE net024 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net024 D VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP13 BEN BE VDD VDD pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 QI_MS QIN_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP3 QI CNN net27 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MP2 net27 QIN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP10 net36 MXI_OUT VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP11 QIN_MS CNN net36 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net32 QI_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 QIN_MS CN net32 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 QIN QI VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP12 CNN CN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP9 QI CN net19 VDD pmos m=1 w=990.00n l=130.00n ng=1 nrd=0 nrs=0
MP8 net19 QI_MS VDD VDD pmos m=1 w=990.00n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWREG4 ACLK_N_I ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX1 A Z VDD VSS
MN1 net010 net032 VSS VSS nmos m=1 w=300.0n l=160.00n ng=1 
+ nrd=0 nrs=0
MN2 net032 A net014 VSS nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MN0 Z net032 net010 VSS nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MN3 net014 A VSS VSS nmos m=1 w=300.0n l=160.00n ng=1 nrd=0 
+ nrs=0
MP1 Z net032 net07 VDD pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
MP3 net011 A VDD VDD pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
MP0 net07 net032 VDD VDD pmos m=1 w=720.00n l=160.00n ng=1 
+ nrd=0 nrs=0
MP2 net032 A net011 VDD pmos m=1 w=720.00n l=160.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX1_DUMMY A Z VDD VSS
MN0 vss_r vdd_r VSS VSS nmos m=1 w=2.49u l=300.0n ng=3 nrd=0 
+ nrs=0
MP0 vdd_r vss_r VDD VDD pmos m=1 w=3.24u l=640.00n ng=2 nrd=0 
+ nrs=0
R0 Z A lvsres w=2.6e-07 l=6e-07
.ENDS

.SUBCKT RSC_IHPSG13_MX2IX1 A0 A1 S ZN VDD VSS
MP4 SN S VDD VDD pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 nrs=0
MP3 ZN SN net12 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 nrs=0
MP2 net12 A1 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 ZN S net17 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 net17 A0 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 SN S VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN3 net13 A1 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 ZN S net13 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net15 A0 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 ZN SN net15 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_DLY_MUX A SEL Z VDD VSS
XI11 net4 Z VDD VSS / RSC_IHPSG13_CINVX2
XI8 A D<3> SEL net4 VDD VSS / RSC_IHPSG13_MX2IX1
XI20<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1
.ENDS
.SUBCKT RSC_IHPSG13_DFNQX2 CN D Q VDD VSS
MN0 Q QIN_SL VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN10 QIN_SL CNN net21 VSS nmos m=1 w=850.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN11 net21 QI_MS VSS VSS nmos m=1 w=850.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN7 net30 QI_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN6 QIN_MS CNN net30 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 QI_MS QIN_MS VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN12 CNN CN VSS VSS nmos m=1 w=495.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN9 net37 D VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN8 QIN_MS CN net37 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 QIN_SL CN net25 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net25 QI_SL VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN2 QI_SL QIN_SL VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP0 Q QIN_SL VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 QI_MS QIN_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP3 QIN_SL CNN net27 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net27 QI_SL VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP10 net36 D VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP11 QIN_MS CNN net36 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net32 QI_MS VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 QIN_MS CN net32 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 QI_SL QIN_SL VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP12 CNN CN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP9 QIN_SL CN net19 VDD pmos m=1 w=990.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP8 net19 QI_MS VDD VDD pmos m=1 w=990.00n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CNAND2X2 A B Z VDD VSS
MN0 Z B net6 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 net6 A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 Z B VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CGATEPX4 CP E Q VDD VSS
MN1 net08 QIN VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net019 net08 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN3 QIN CP net019 VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 nrs=0
MN6 Q net015 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 
+ nrs=0
MN5 net015 net08 net018 VSS nmos m=1 w=980.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MN8 QIN CPN net023 VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN7 net023 E VSS VSS nmos m=1 w=870.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net018 CP VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 CPN CP VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP3 net08 QIN VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 QIN CPN net017 VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net017 net08 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 
+ nrd=0 nrs=0
MP0 CPN CP VDD VDD pmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP8 QIN CP net024 VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 net024 E VDD VDD pmos m=1 w=975.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net015 CP VDD VDD pmos m=1 w=1.27u l=130.00n ng=1 nrd=0 
+ nrs=0
MP6 Q net015 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 
+ nrs=0
MP5 net015 net08 VDD VDD pmos m=1 w=1.27u l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CBUFX8 A Z VDD VSS
MP0 net4 A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net4 VDD VDD pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
MN1 Z net4 VSS VSS nmos m=1 w=2.82u l=130.00n ng=4 nrd=0 nrs=0
MN0 net4 A VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CDLYX2 A Z VDD VSS
MN2 net4 A net9 VSS nmos m=1 w=320.00n l=200.0n ng=1 nrd=0 nrs=0
MN0 Z net4 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net9 A VSS VSS nmos m=1 w=320.00n l=200.0n ng=1 nrd=0 nrs=0
MP2 net4 A net10 VDD pmos m=1 w=1.2u l=200.0n ng=1 nrd=0 nrs=0
MP1 net10 A VDD VDD pmos m=1 w=1.2u l=200.0n ng=1 nrd=0 nrs=0
MP0 Z net4 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MX2X2 A0 A1 S Z VDD VSS
MP6 Z net010 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 SN S VDD VDD pmos m=1 w=645.000n l=130.00n ng=1 nrd=0 nrs=0
MP3 net010 SN net12 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net12 A1 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net010 S net17 VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net17 A0 VDD VDD pmos m=1 w=985.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 Z net010 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 SN S VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 nrs=0
MN3 net13 A1 VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net010 S net13 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net15 A0 VSS VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net010 SN net15 VSS nmos m=1 w=560.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_AND2X2 A B Z VDD VSS
MN3 Z net6 VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net9 B VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net6 B VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_TIEL Z VDD VSS
MN0 Z net2 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 net2 net2 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_XOR2X2 A B Z VDD VSS
MP8 net012 B net7 VDD pmos m=1 w=825.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP7 net011 net3 net012 VDD pmos m=1 w=825.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP6 Z net012 VDD VDD pmos m=1 w=1.535u l=130.00n ng=1 nrd=0 
+ nrs=0
MP2 net7 A VDD VDD pmos m=1 w=825.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP4 net011 net7 VDD VDD pmos m=1 w=825.000n l=130.00n ng=1 
+ nrd=0 nrs=0
MP5 net3 B VDD VDD pmos m=1 w=580.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN7 net012 B net011 VSS nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN6 net7 net3 net012 VSS nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN5 Z net012 VSS VSS nmos m=1 w=775.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN2 net7 A VSS VSS nmos m=1 w=555.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN4 net3 B VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 net011 net7 VSS VSS nmos m=1 w=555.000n l=130.00n ng=1 
+ nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_OA12X1 A B C Z VDD VSS
MN2 net7 C VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN3 Z net17 VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MN1 net17 B net7 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN0 net17 A net7 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 net24 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP3 Z net17 VDD VDD pmos m=1 w=905.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net17 B net24 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP2 net17 C VDD VDD pmos m=1 w=905.000n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_CTRL ACLK_N BIST_CK_I BIST_CS_I BIST_EN BIST_RE_I 
+ BIST_WE_I B_TIEL_O CK_I CS_I DCLK ECLK PULSE_H PULSE_L PULSE_O RCLK RE_I 
+ ROW_CS WCLK WE_I VDD VSS
XI17 ck_regs we col_we VDD VSS / RSC_IHPSG13_DFNQX2
XI16 ck_regs re col_re VDD VSS / RSC_IHPSG13_DFNQX2
XI18 ck_regs cs net7 VDD VSS / RSC_IHPSG13_DFNQX2
XI71 ACLK_N net012 PULSE_O VDD VSS / RSC_IHPSG13_DFNQX2
XI77 col_we net9 net016 VDD VSS / RSC_IHPSG13_CNAND2X2
XI76 col_re net9 net018 VDD VSS / RSC_IHPSG13_CNAND2X2
XI15 ck_dly WEorREandCS aclk VDD VSS / RSC_IHPSG13_CGATEPX4
XI14 ck WEandCS DCLK VDD VSS / RSC_IHPSG13_CGATEPX4
XI60 net7 ROW_CS VDD VSS / RSC_IHPSG13_CBUFX8
XI73 PULSE_O net012 VDD VSS / RSC_IHPSG13_CINVX2
XI8 net9 net8 VDD VSS / RSC_IHPSG13_CINVX2
XI64 ck ck_dly VDD VSS / RSC_IHPSG13_CDLYX2
XI86 CS_I BIST_CS_I BIST_EN cs VDD VSS / RSC_IHPSG13_MX2X2
XI87 CK_I BIST_CK_I BIST_EN ck VDD VSS / RSC_IHPSG13_MX2X2
XI85 WE_I BIST_WE_I BIST_EN we VDD VSS / RSC_IHPSG13_MX2X2
XI84 RE_I BIST_RE_I BIST_EN re VDD VSS / RSC_IHPSG13_MX2X2
XI22 we cs WEandCS VDD VSS / RSC_IHPSG13_AND2X2
XBM_TIEL B_TIEL_O VDD VSS / RSC_IHPSG13_TIEL
XI48 ck_dly ck_regs VDD VSS / RSC_IHPSG13_CINVX4
XI81 net016 WCLK VDD VSS / RSC_IHPSG13_CINVX4
XI80 net018 RCLK VDD VSS / RSC_IHPSG13_CINVX4
XI78 net8 net020 VDD VSS / RSC_IHPSG13_CINVX4
XI6 PULSE_L PULSE_H net9 VDD VSS / RSC_IHPSG13_XOR2X2
XI79 net020 ECLK VDD VSS / RSC_IHPSG13_CINVX8
XI63 aclk ACLK_N VDD VSS / RSC_IHPSG13_CINVX8
XI21 re we cs WEorREandCS VDD VSS / RSC_IHPSG13_OA12X1
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDEC2 ACLK_N ADDR<1> ADDR<0> ADDR_COL<1> ADDR_COL<0> 
+ ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> ADDR_DEC<2> 
+ ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI14<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI14<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net6<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net6<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<3> PADR<1> PADR<0> addr_n<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<2> PADR<1> NADR<0> addr_n<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<1> NADR<1> PADR<0> addr_n<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<0> NADR<1> NADR<0> addr_n<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI16<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI17<3> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_TIEL
XI17<2> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_TIEL
XI17<1> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_TIEL
XI17<0> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RSC_IHPSG13_NOR2X2 A B Z VDD VSS
MP1 Z B net9 VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net9 A VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MN0 Z B VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN1 Z A VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CINVX4_WN A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BLDRV BLC BLC_SEL BLT BLT_SEL PRE_N SEL_P WR_ONE WR_ZERO 
+ VDD VSS
XCDEC SEL_P WR_ZERO BLC_PMOS_DRIVE VDD VSS / RSC_IHPSG13_NAND2X2
XTDEC SEL_P WR_ONE BLT_PMOS_DRIVE VDD VSS / RSC_IHPSG13_NAND2X2
MTWN BLT BLT_NMOS_DRIVE VSS VSS nmos m=1 w=4.82u l=130.00n 
+ ng=2 nrd=0 nrs=0
MCWN BLC BLC_NMOS_DRIVE VSS VSS nmos m=1 w=4.82u l=130.00n 
+ ng=2 nrd=0 nrs=0
MCWP BLC BLC_PMOS_DRIVE VDD VDD pmos m=1 w=1.5u l=130.00n ng=1 
+ nrd=0 nrs=0
MTWP BLT BLT_PMOS_DRIVE VDD VDD pmos m=1 w=1.5u l=130.00n ng=1 
+ nrd=0 nrs=0
MTSP BLT_SEL SEL_N BLT VDD pmos m=1 w=1.5u l=130.00n ng=1 nrd=0 
+ nrs=0
MTPR BLT PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n ng=2 nrd=0 
+ nrs=0
MCSP BLC_SEL SEL_N BLC VDD pmos m=1 w=1.5u l=130.00n ng=1 nrd=0 
+ nrs=0
MCPR BLC PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n ng=2 nrd=0 
+ nrs=0
XI86 SEL_P SEL_N VDD VSS / RSC_IHPSG13_INVX2
XTINV BLC_PMOS_DRIVE BLT_NMOS_DRIVE VDD VSS / RSC_IHPSG13_INVX2
XCINV BLT_PMOS_DRIVE BLC_NMOS_DRIVE VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RSC_IHPSG13_TIEH Z VDD VSS
MN0 net2 net2 VSS VSS nmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP0 Z net2 VDD VDD pmos m=1 w=480.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_MET3RES A B
R0 B A lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RSC_IHPSG13_DFPQD_MSAFFX2 CP DN DP QN QP VDD VSS
MN12 SN RN DIFFP VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN13 TAIL CP VSS VSS nmos m=1 w=2.4u l=130.00n ng=2 nrd=0 nrs=0
MN9 DIFFP DP TAIL VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN10 DIFFN DN TAIL VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN11 RN SN DIFFN VSS nmos m=1 w=2.4u l=200.0n ng=2 nrd=0 nrs=0
MN19 net33 SN VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN20 QN QP net37 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MN18 net37 RN VSS VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MN17 QP QN net33 VSS nmos m=1 w=980.00n l=130.00n ng=1 nrd=0 nrs=0
MP15 SN RN VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP16 RN CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP14 DIFFP CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MP12 RN SN VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP13 DIFFN CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 
+ nrs=0
MP11 SN CP VDD VDD pmos m=1 w=800.0n l=130.00n ng=1 nrd=0 nrs=0
MP19 QN QP VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
MP20 QP SN VDD VDD pmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP18 QN RN VDD VDD pmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP17 QP QN VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_CBUFX2 A Z VDD VSS
MN1 Z net4 VSS VSS nmos m=1 w=705.000n l=130.00n ng=1 nrd=0 
+ nrs=0
MN0 net4 A VSS VSS nmos m=1 w=540.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 Z net4 VDD VDD pmos m=1 w=1.62u l=130.00n ng=1 nrd=0 nrs=0
MP0 net4 A VDD VDD pmos m=1 w=1.1u l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RSC_IHPSG13_INVX4 A Z VDD VSS
MN0 Z A VSS VSS nmos m=1 w=1.96u l=130.00n ng=2 nrd=0 nrs=0
MP0 Z A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLCTRL2 A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<3> A_BLC<2> A_BLC<1> 
+ A_BLC<0> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I80 A_WCLK_B_R A_RCLK_B_R net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I44 A_WCLK_B_R A_BM_N A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_ADDR_DEC<2> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_ADDR_DEC<1> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<0> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_R A_RCLK_B_L / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_R A_RCLK_L / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_R A_WCLK_B_L / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I78 A_RCLK_B_R A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_R VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_R A_RCLK_B_R VDD VSS / RSC_IHPSG13_CINVX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4 VDD VSS
XI0<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2 VDD VSS
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDEC4 ACLK_N ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<3> BIST_ADDR<2> 
+ BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI15 ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI14 addr_int ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int net7<0> VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RSC_IHPSG13_AND2X4 A B Z VDD VSS
MN3 Z net6 VSS VSS nmos m=1 w=1.96u l=130.00n ng=2 nrd=0 nrs=0
MN4 net9 B VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
MP0 net6 B VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLCTRL4 A_ADDR_COL A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<15> A_BLC<14> 
+ A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> 
+ A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> 
+ A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L 
+ A_DCLK_B_R A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L 
+ A_RCLK_R A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_I80 A_WCLK_B_L A_RCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DO_WRITE_P A_DI_N A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XA_CAPS<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_N0 A_P0 VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL A_N0 VDD VSS / RSC_IHPSG13_CINVX4
XA_I81<1> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<15> A_BLC<15> A_BLC_SEL A_BLT<15> A_BLT_SEL A_PRE_N A_SEL_P<15> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<14> A_BLC<14> A_BLC_SEL A_BLT<14> A_BLT_SEL A_PRE_N A_SEL_P<14> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<13> A_BLC<13> A_BLC_SEL A_BLT<13> A_BLT_SEL A_PRE_N A_SEL_P<13> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<12> A_BLC<12> A_BLC_SEL A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<12> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<11> A_BLC<11> A_BLC_SEL A_BLT<11> A_BLT_SEL A_PRE_N A_SEL_P<11> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<10> A_BLC<10> A_BLC_SEL A_BLT<10> A_BLT_SEL A_PRE_N A_SEL_P<10> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<9> A_BLC<9> A_BLC_SEL A_BLT<9> A_BLT_SEL A_PRE_N A_SEL_P<9> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<8> A_BLC<8> A_BLC_SEL A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<8> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_SEL_P<7> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_SEL_P<6> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_SEL_P<5> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<4> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_SEL_P<3> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_SEL_P<2> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_SEL_P<1> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<0> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net24 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3INV<15> net23<0> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<1> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<2> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<3> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<4> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<5> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<6> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<7> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<8> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<9> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<10> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<11> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<12> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<13> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<14> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<15> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I70<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI73<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_DEC3<15> A_P0 A_ADDR_DEC<7> net23<0> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<14> A_P0 A_ADDR_DEC<6> net23<1> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<13> A_P0 A_ADDR_DEC<5> net23<2> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<12> A_P0 A_ADDR_DEC<4> net23<3> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<11> A_P0 A_ADDR_DEC<3> net23<4> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<10> A_P0 A_ADDR_DEC<2> net23<5> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<9> A_P0 A_ADDR_DEC<1> net23<6> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<8> A_P0 A_ADDR_DEC<0> net23<7> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<7> A_N0 A_ADDR_DEC<7> net23<8> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<6> A_N0 A_ADDR_DEC<6> net23<9> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<5> A_N0 A_ADDR_DEC<5> net23<10> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<4> A_N0 A_ADDR_DEC<4> net23<11> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<3> A_N0 A_ADDR_DEC<3> net23<12> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<2> A_N0 A_ADDR_DEC<2> net23<13> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<1> A_N0 A_ADDR_DEC<1> net23<14> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<0> A_N0 A_ADDR_DEC<0> net23<15> VDD VSS / RSC_IHPSG13_NAND2X2
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDEC3 ACLK_N ADDR<2> ADDR<1> ADDR<0> ADDR_COL<1> 
+ ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> 
+ ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> 
+ BIST_EN_I VDD VSS
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net6<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net6<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net6<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLCTRL3 A_ADDR_DEC<7> A_ADDR_DEC<6> A_ADDR_DEC<5> 
+ A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> A_ADDR_DEC<0> 
+ A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> 
+ A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R A_DCLK_L 
+ A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R A_TIEH_O 
+ A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_R A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_I70<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I70<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I44 A_BM_N A_WCLK_B_R A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_ADDR_DEC<7> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_ADDR_DEC<6> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_ADDR_DEC<5> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_ADDR_DEC<4> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_ADDR_DEC<2> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_ADDR_DEC<1> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<0> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I80 A_WCLK_B_R A_RCLK_B_R net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_16x2_CORNER VDD_CORE VSS
XI16 VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR A_WL B_WL NW PW VDD VSS
MN1 VSS A_WL VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 VSS B_WL VSS VSS nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_16x2_EDGE_LR A_WL<15> A_WL<14> A_WL<13> A_WL<12> 
+ A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> 
+ A_WL<2> A_WL<1> A_WL<0> B_WL<15> B_WL<14> B_WL<13> B_WL<12> B_WL<11> 
+ B_WL<10> B_WL<9> B_WL<8> B_WL<7> B_WL<6> B_WL<5> B_WL<4> B_WL<3> B_WL<2> 
+ B_WL<1> B_WL<0> VDD_CORE VSS
XI0<15> A_WL<15> B_WL<15> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<14> A_WL<14> B_WL<14> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<13> A_WL<13> B_WL<13> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<12> A_WL<12> B_WL<12> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<11> A_WL<11> B_WL<11> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<10> A_WL<10> B_WL<10> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<9> A_WL<9> B_WL<9> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<8> A_WL<8> B_WL<8> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<7> A_WL<7> B_WL<7> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<6> A_WL<6> B_WL<6> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<5> A_WL<5> B_WL<5> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<4> A_WL<4> B_WL<4> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<3> A_WL<3> B_WL<3> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<2> A_WL<2> B_WL<2> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<1> A_WL<1> B_WL<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
XI0<0> A_WL<0> B_WL<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_LR
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL A_BLC_BOT A_BLC_TOP A_BLT_BOT A_BLT_TOP 
+ A_LWL A_RWL B_BLC_BOT B_BLC_TOP B_BLT_BOT B_BLT_TOP B_LWL B_RWL NW PW VDD VSS
MN5 NC B_RWL B_BLC_BOT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN4 B_BLT_BOT B_LWL NT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN0 NC NT VSS PW nmos m=1 w=600.0n l=130.00n ng=2 nrd=0 nrs=0
MN1 NT NC VSS PW nmos m=1 w=600.0n l=130.00n ng=2 nrd=0 nrs=0
MN3 NC A_RWL A_BLC_TOP PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MN2 A_BLT_TOP A_LWL NT PW nmos m=1 w=300.0n l=130.00n ng=1 nrd=0 nrs=0
MP1 NT NC VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
MP0 NC NT VDD NW pmos m=1 w=150.00n l=130.00n ng=1 nrd=0 nrs=0
R5 B_RWL B_LWL lvsres w=2.6e-07 l=6e-07
R4 B_BLC_BOT B_BLC_TOP lvsres w=2.6e-07 l=6e-07
R3 B_BLT_BOT B_BLT_TOP lvsres w=2.6e-07 l=6e-07
R1 A_BLC_BOT A_BLC_TOP lvsres w=2.6e-07 l=6e-07
R0 A_BLT_BOT A_BLT_TOP lvsres w=2.6e-07 l=6e-07
R2 A_RWL A_LWL lvsres w=2.6e-07 l=6e-07
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_16x2_SRAM A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> 
+ A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<15> 
+ A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> 
+ A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> 
+ A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> 
+ A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> B_BLC_BOT<1> 
+ B_BLC_BOT<0> B_BLC_TOP<1> B_BLC_TOP<0> B_BLT_BOT<1> B_BLT_BOT<0> 
+ B_BLT_TOP<1> B_BLT_TOP<0> B_LWL<15> B_LWL<14> B_LWL<13> B_LWL<12> B_LWL<11> 
+ B_LWL<10> B_LWL<9> B_LWL<8> B_LWL<7> B_LWL<6> B_LWL<5> B_LWL<4> B_LWL<3> 
+ B_LWL<2> B_LWL<1> B_LWL<0> B_RWL<15> B_RWL<14> B_RWL<13> B_RWL<12> B_RWL<11> 
+ B_RWL<10> B_RWL<9> B_RWL<8> B_RWL<7> B_RWL<6> B_RWL<5> B_RWL<4> B_RWL<3> 
+ B_RWL<2> B_RWL<1> B_RWL<0> VDD_CORE VSS
XCELL<31> A_BLC_TOP<1> A_RBLC<15> A_BLT_TOP<1> A_RBLT<15> A_XWL<15> A_RWL<15> 
+ B_BLC_TOP<1> B_RBLC<15> B_BLT_TOP<1> B_RBLT<15> B_XWL<15> B_RWL<15> 
+ VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<30> A_RBLC<14> A_RBLC<15> A_RBLT<14> A_RBLT<15> A_XWL<14> A_RWL<14> 
+ B_RBLC<14> B_RBLC<15> B_RBLT<14> B_RBLT<15> B_XWL<14> B_RWL<14> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<29> A_RBLC<14> A_RBLC<13> A_RBLT<14> A_RBLT<13> A_XWL<13> A_RWL<13> 
+ B_RBLC<14> B_RBLC<13> B_RBLT<14> B_RBLT<13> B_XWL<13> B_RWL<13> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<28> A_RBLC<12> A_RBLC<13> A_RBLT<12> A_RBLT<13> A_XWL<12> A_RWL<12> 
+ B_RBLC<12> B_RBLC<13> B_RBLT<12> B_RBLT<13> B_XWL<12> B_RWL<12> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<27> A_RBLC<12> A_RBLC<11> A_RBLT<12> A_RBLT<11> A_XWL<11> A_RWL<11> 
+ B_RBLC<12> B_RBLC<11> B_RBLT<12> B_RBLT<11> B_XWL<11> B_RWL<11> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<26> A_RBLC<10> A_RBLC<11> A_RBLT<10> A_RBLT<11> A_XWL<10> A_RWL<10> 
+ B_RBLC<10> B_RBLC<11> B_RBLT<10> B_RBLT<11> B_XWL<10> B_RWL<10> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<25> A_RBLC<10> A_RBLC<9> A_RBLT<10> A_RBLT<9> A_XWL<9> A_RWL<9> 
+ B_RBLC<10> B_RBLC<9> B_RBLT<10> B_RBLT<9> B_XWL<9> B_RWL<9> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<24> A_RBLC<8> A_RBLC<9> A_RBLT<8> A_RBLT<9> A_XWL<8> A_RWL<8> B_RBLC<8> 
+ B_RBLC<9> B_RBLT<8> B_RBLT<9> B_XWL<8> B_RWL<8> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<23> A_RBLC<8> A_RBLC<7> A_RBLT<8> A_RBLT<7> A_XWL<7> A_RWL<7> B_RBLC<8> 
+ B_RBLC<7> B_RBLT<8> B_RBLT<7> B_XWL<7> B_RWL<7> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<22> A_RBLC<6> A_RBLC<7> A_RBLT<6> A_RBLT<7> A_XWL<6> A_RWL<6> B_RBLC<6> 
+ B_RBLC<7> B_RBLT<6> B_RBLT<7> B_XWL<6> B_RWL<6> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<21> A_RBLC<6> A_RBLC<5> A_RBLT<6> A_RBLT<5> A_XWL<5> A_RWL<5> B_RBLC<6> 
+ B_RBLC<5> B_RBLT<6> B_RBLT<5> B_XWL<5> B_RWL<5> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<20> A_RBLC<4> A_RBLC<5> A_RBLT<4> A_RBLT<5> A_XWL<4> A_RWL<4> B_RBLC<4> 
+ B_RBLC<5> B_RBLT<4> B_RBLT<5> B_XWL<4> B_RWL<4> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<19> A_RBLC<4> A_RBLC<3> A_RBLT<4> A_RBLT<3> A_XWL<3> A_RWL<3> B_RBLC<4> 
+ B_RBLC<3> B_RBLT<4> B_RBLT<3> B_XWL<3> B_RWL<3> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<18> A_RBLC<2> A_RBLC<3> A_RBLT<2> A_RBLT<3> A_XWL<2> A_RWL<2> B_RBLC<2> 
+ B_RBLC<3> B_RBLT<2> B_RBLT<3> B_XWL<2> B_RWL<2> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<17> A_RBLC<2> A_RBLC<1> A_RBLT<2> A_RBLT<1> A_XWL<1> A_RWL<1> B_RBLC<2> 
+ B_RBLC<1> B_RBLT<2> B_RBLT<1> B_XWL<1> B_RWL<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<16> A_BLC_BOT<1> A_RBLC<1> A_BLT_BOT<1> A_RBLT<1> A_XWL<0> A_RWL<0> 
+ B_BLC_BOT<1> B_RBLC<1> B_BLT_BOT<1> B_RBLT<1> B_XWL<0> B_RWL<0> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<15> A_BLC_TOP<0> A_LBLC<15> A_BLT_TOP<0> A_LBLT<15> A_LWL<15> A_XWL<15> 
+ B_BLC_TOP<0> B_LBLC<15> B_BLT_TOP<0> B_LBLT<15> B_LWL<15> B_XWL<15> 
+ VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<14> A_LBLC<14> A_LBLC<15> A_LBLT<14> A_LBLT<15> A_LWL<14> A_XWL<14> 
+ B_LBLC<14> B_LBLC<15> B_LBLT<14> B_LBLT<15> B_LWL<14> B_XWL<14> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<13> A_LBLC<14> A_LBLC<13> A_LBLT<14> A_LBLT<13> A_LWL<13> A_XWL<13> 
+ B_LBLC<14> B_LBLC<13> B_LBLT<14> B_LBLT<13> B_LWL<13> B_XWL<13> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<12> A_LBLC<12> A_LBLC<13> A_LBLT<12> A_LBLT<13> A_LWL<12> A_XWL<12> 
+ B_LBLC<12> B_LBLC<13> B_LBLT<12> B_LBLT<13> B_LWL<12> B_XWL<12> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<11> A_LBLC<12> A_LBLC<11> A_LBLT<12> A_LBLT<11> A_LWL<11> A_XWL<11> 
+ B_LBLC<12> B_LBLC<11> B_LBLT<12> B_LBLT<11> B_LWL<11> B_XWL<11> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<10> A_LBLC<10> A_LBLC<11> A_LBLT<10> A_LBLT<11> A_LWL<10> A_XWL<10> 
+ B_LBLC<10> B_LBLC<11> B_LBLT<10> B_LBLT<11> B_LWL<10> B_XWL<10> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<9> A_LBLC<10> A_LBLC<9> A_LBLT<10> A_LBLT<9> A_LWL<9> A_XWL<9> 
+ B_LBLC<10> B_LBLC<9> B_LBLT<10> B_LBLT<9> B_LWL<9> B_XWL<9> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<8> A_LBLC<8> A_LBLC<9> A_LBLT<8> A_LBLT<9> A_LWL<8> A_XWL<8> B_LBLC<8> 
+ B_LBLC<9> B_LBLT<8> B_LBLT<9> B_LWL<8> B_XWL<8> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<7> A_LBLC<8> A_LBLC<7> A_LBLT<8> A_LBLT<7> A_LWL<7> A_XWL<7> B_LBLC<8> 
+ B_LBLC<7> B_LBLT<8> B_LBLT<7> B_LWL<7> B_XWL<7> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<6> A_LBLC<6> A_LBLC<7> A_LBLT<6> A_LBLT<7> A_LWL<6> A_XWL<6> B_LBLC<6> 
+ B_LBLC<7> B_LBLT<6> B_LBLT<7> B_LWL<6> B_XWL<6> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<5> A_LBLC<6> A_LBLC<5> A_LBLT<6> A_LBLT<5> A_LWL<5> A_XWL<5> B_LBLC<6> 
+ B_LBLC<5> B_LBLT<6> B_LBLT<5> B_LWL<5> B_XWL<5> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<4> A_LBLC<4> A_LBLC<5> A_LBLT<4> A_LBLT<5> A_LWL<4> A_XWL<4> B_LBLC<4> 
+ B_LBLC<5> B_LBLT<4> B_LBLT<5> B_LWL<4> B_XWL<4> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<3> A_LBLC<4> A_LBLC<3> A_LBLT<4> A_LBLT<3> A_LWL<3> A_XWL<3> B_LBLC<4> 
+ B_LBLC<3> B_LBLT<4> B_LBLT<3> B_LWL<3> B_XWL<3> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<2> A_LBLC<2> A_LBLC<3> A_LBLT<2> A_LBLT<3> A_LWL<2> A_XWL<2> B_LBLC<2> 
+ B_LBLC<3> B_LBLT<2> B_LBLT<3> B_LWL<2> B_XWL<2> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<1> A_LBLC<2> A_LBLC<1> A_LBLT<2> A_LBLT<1> A_LWL<1> A_XWL<1> B_LBLC<2> 
+ B_LBLC<1> B_LBLT<2> B_LBLT<1> B_LWL<1> B_XWL<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
XCELL<0> A_BLC_BOT<0> A_LBLC<1> A_BLT_BOT<0> A_LBLT<1> A_LWL<0> A_XWL<0> 
+ B_BLC_BOT<0> B_LBLC<1> B_BLT_BOT<0> B_LBLT<1> B_LWL<0> B_XWL<0> VDD_CORE 
+ VSS VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_CELL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB A_BLC A_BLT B_BLC B_BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_16x2_EDGE_TB A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ B_BLC<1> B_BLC<0> B_BLT<1> B_BLT<0> VDD_CORE VSS
XEDGE<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB
XEDGE<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_TAP A_BLC A_BLT B_BLC B_BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_16x2_TAP A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ B_BLC<1> B_BLC<0> B_BLT<1> B_BLT<0> VDD_CORE VSS
XIEDGEBP_COL1<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL1<0> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL2<1> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB
XIEDGEBP_COL2<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_EDGE_TB
XITAP<1> A_BLC<1> A_BLT<1> B_BLC<1> B_BLT<1> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_TAP
XITAP<0> A_BLC<0> A_BLT<0> B_BLC<0> B_BLT<0> VDD_CORE VSS 
+ VDD_CORE VSS / RM_IHPSG13_2048x64_c2_2P_BITKIT_TAP
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_TAP_LR NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BITKIT_16x2_TAP_LR VDD_CORE VSS
XCORNER<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER
XCORNER<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER
XTAP_BORDER VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_TAP_LR
.ENDS

.SUBCKT RSC_IHPSG13_CBUFX12 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=4.23u l=130.00n ng=6 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=9.72u l=130.00n ng=6 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=3.24u l=130.00n ng=2 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDRV13X12 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX12 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=9.72u l=130.00n ng=6 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_WLDRV16X12 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX12
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_DEC04 ADDR<3> ADDR<2> ADDR<1> ADDR<0> CS ECLK_H_BOT 
+ ECLK_H_TOP ECLK_L_BOT ECLK_L_TOP WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> 
+ WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> VDD VSS
XI0<3> PADR<1> PADR<0> sel01<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<2> PADR<1> NADR<0> sel01<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<1> NADR<1> PADR<0> sel01<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI0<0> NADR<1> NADR<0> sel01<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI4 ECLK_L_BOT EN VDD VSS / RSC_IHPSG13_CINVX4
XI5 ECLK_H_BOT ECLK_L_BOT VDD VSS / RSC_IHPSG13_CINVX2
XI3<3> PADR<3> NADR<3> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> PADR<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> PADR<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> PADR<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XR0 ECLK_H_BOT ECLK_H_TOP / RSC_IHPSG13_MET2RES
XI11 ECLK_L_BOT ECLK_L_TOP / RSC_IHPSG13_MET2RES
XI1<3> PADR<2> PADR<3> CS sel23<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<2> PADR<3> CS sel23<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<2> NADR<3> CS sel23<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<2> NADR<3> CS sel23<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI2<15> sel23<3> sel01<3> EN WL<15> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<14> sel23<3> sel01<2> EN WL<14> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<13> sel23<3> sel01<1> EN WL<13> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<12> sel23<3> sel01<0> EN WL<12> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<11> sel23<2> sel01<3> EN WL<11> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<10> sel23<2> sel01<2> EN WL<10> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<9> sel23<2> sel01<1> EN WL<9> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<8> sel23<2> sel01<0> EN WL<8> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<7> sel23<1> sel01<3> EN WL<7> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<6> sel23<1> sel01<2> EN WL<6> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<5> sel23<1> sel01<1> EN WL<5> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<4> sel23<1> sel01<0> EN WL<4> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<3> sel23<0> sel01<3> EN WL<3> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<2> sel23<0> sel01<2> EN WL<2> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<1> sel23<0> sel01<1> EN WL<1> VDD VSS / RSC_IHPSG13_NOR3X2
XI2<0> sel23<0> sel01<0> EN WL<0> VDD VSS / RSC_IHPSG13_NOR3X2
XCAPS4 VDD VSS / RSC_IHPSG13_FILLCAP4
XLATCH<3> CS ADDR<3> PADR<3> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<2> CS ADDR<2> PADR<2> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<1> CS ADDR<1> PADR<1> VDD VSS / RSC_IHPSG13_LHPQX2
XLATCH<0> CS ADDR<0> PADR<0> VDD VSS / RSC_IHPSG13_LHPQX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_DEC02 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC ADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI2<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI2<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_DEC01 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC NADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI2<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI2<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_DEC00 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC NADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV<1> ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XADDRINV<0> ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_DEC03 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDEC ADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWDEC9 ADDR_N_I<8> ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> 
+ ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I 
+ WL_O<511> WL_O<510> WL_O<509> WL_O<508> WL_O<507> WL_O<506> WL_O<505> 
+ WL_O<504> WL_O<503> WL_O<502> WL_O<501> WL_O<500> WL_O<499> WL_O<498> 
+ WL_O<497> WL_O<496> WL_O<495> WL_O<494> WL_O<493> WL_O<492> WL_O<491> 
+ WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> WL_O<484> 
+ WL_O<483> WL_O<482> WL_O<481> WL_O<480> WL_O<479> WL_O<478> WL_O<477> 
+ WL_O<476> WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> 
+ WL_O<469> WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> WL_O<463> 
+ WL_O<462> WL_O<461> WL_O<460> WL_O<459> WL_O<458> WL_O<457> WL_O<456> 
+ WL_O<455> WL_O<454> WL_O<453> WL_O<452> WL_O<451> WL_O<450> WL_O<449> 
+ WL_O<448> WL_O<447> WL_O<446> WL_O<445> WL_O<444> WL_O<443> WL_O<442> 
+ WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> WL_O<436> WL_O<435> 
+ WL_O<434> WL_O<433> WL_O<432> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> WL_O<415> WL_O<414> 
+ WL_O<413> WL_O<412> WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> 
+ WL_O<406> WL_O<405> WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> 
+ WL_O<399> WL_O<398> WL_O<397> WL_O<396> WL_O<395> WL_O<394> WL_O<393> 
+ WL_O<392> WL_O<391> WL_O<390> WL_O<389> WL_O<388> WL_O<387> WL_O<386> 
+ WL_O<385> WL_O<384> WL_O<383> WL_O<382> WL_O<381> WL_O<380> WL_O<379> 
+ WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> WL_O<372> 
+ WL_O<371> WL_O<370> WL_O<369> WL_O<368> WL_O<367> WL_O<366> WL_O<365> 
+ WL_O<364> WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> 
+ WL_O<357> WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> WL_O<351> 
+ WL_O<350> WL_O<349> WL_O<348> WL_O<347> WL_O<346> WL_O<345> WL_O<344> 
+ WL_O<343> WL_O<342> WL_O<341> WL_O<340> WL_O<339> WL_O<338> WL_O<337> 
+ WL_O<336> WL_O<335> WL_O<334> WL_O<333> WL_O<332> WL_O<331> WL_O<330> 
+ WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> WL_O<324> WL_O<323> 
+ WL_O<322> WL_O<321> WL_O<320> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> WL_O<303> WL_O<302> 
+ WL_O<301> WL_O<300> WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> 
+ WL_O<294> WL_O<293> WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> 
+ WL_O<287> WL_O<286> WL_O<285> WL_O<284> WL_O<283> WL_O<282> WL_O<281> 
+ WL_O<280> WL_O<279> WL_O<278> WL_O<277> WL_O<276> WL_O<275> WL_O<274> 
+ WL_O<273> WL_O<272> WL_O<271> WL_O<270> WL_O<269> WL_O<268> WL_O<267> 
+ WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> WL_O<260> 
+ WL_O<259> WL_O<258> WL_O<257> WL_O<256> WL_O<255> WL_O<254> WL_O<253> 
+ WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> 
+ WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> WL_O<239> 
+ WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> WL_O<233> WL_O<232> 
+ WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> WL_O<226> WL_O<225> 
+ WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> WL_O<219> WL_O<218> 
+ WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> WL_O<212> WL_O<211> 
+ WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> WL_O<191> WL_O<190> 
+ WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> 
+ WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> 
+ WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> WL_O<170> WL_O<169> 
+ WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> WL_O<163> WL_O<162> 
+ WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> WL_O<156> WL_O<155> 
+ WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> WL_O<148> 
+ WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> WL_O<142> WL_O<141> 
+ WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> 
+ WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> WL_O<127> 
+ WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> 
+ WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> 
+ WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> 
+ WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> 
+ WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XSEL<31> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<31> ECLK_H<31> 
+ ECLK_H<32> ECLK_B<31> ECLK_B<32> WL_O<511> WL_O<510> WL_O<509> WL_O<508> 
+ WL_O<507> WL_O<506> WL_O<505> WL_O<504> WL_O<503> WL_O<502> WL_O<501> 
+ WL_O<500> WL_O<499> WL_O<498> WL_O<497> WL_O<496> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<30> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<30> ECLK_H<30> 
+ ECLK_H<31> ECLK_B<30> ECLK_B<31> WL_O<495> WL_O<494> WL_O<493> WL_O<492> 
+ WL_O<491> WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> 
+ WL_O<484> WL_O<483> WL_O<482> WL_O<481> WL_O<480> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<29> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<29> ECLK_H<29> 
+ ECLK_H<30> ECLK_B<29> ECLK_B<30> WL_O<479> WL_O<478> WL_O<477> WL_O<476> 
+ WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> WL_O<469> 
+ WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<28> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<28> ECLK_H<28> 
+ ECLK_H<29> ECLK_B<28> ECLK_B<29> WL_O<463> WL_O<462> WL_O<461> WL_O<460> 
+ WL_O<459> WL_O<458> WL_O<457> WL_O<456> WL_O<455> WL_O<454> WL_O<453> 
+ WL_O<452> WL_O<451> WL_O<450> WL_O<449> WL_O<448> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<27> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<27> ECLK_H<27> 
+ ECLK_H<28> ECLK_B<27> ECLK_B<28> WL_O<447> WL_O<446> WL_O<445> WL_O<444> 
+ WL_O<443> WL_O<442> WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> 
+ WL_O<436> WL_O<435> WL_O<434> WL_O<433> WL_O<432> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<26> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<26> ECLK_H<26> 
+ ECLK_H<27> ECLK_B<26> ECLK_B<27> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<25> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<25> ECLK_H<25> 
+ ECLK_H<26> ECLK_B<25> ECLK_B<26> WL_O<415> WL_O<414> WL_O<413> WL_O<412> 
+ WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> WL_O<406> WL_O<405> 
+ WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<24> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<24> ECLK_H<24> 
+ ECLK_H<25> ECLK_B<24> ECLK_B<25> WL_O<399> WL_O<398> WL_O<397> WL_O<396> 
+ WL_O<395> WL_O<394> WL_O<393> WL_O<392> WL_O<391> WL_O<390> WL_O<389> 
+ WL_O<388> WL_O<387> WL_O<386> WL_O<385> WL_O<384> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<23> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<23> ECLK_H<23> 
+ ECLK_H<24> ECLK_B<23> ECLK_B<24> WL_O<383> WL_O<382> WL_O<381> WL_O<380> 
+ WL_O<379> WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> 
+ WL_O<372> WL_O<371> WL_O<370> WL_O<369> WL_O<368> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<22> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<22> ECLK_H<22> 
+ ECLK_H<23> ECLK_B<22> ECLK_B<23> WL_O<367> WL_O<366> WL_O<365> WL_O<364> 
+ WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> WL_O<357> 
+ WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<21> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<21> ECLK_H<21> 
+ ECLK_H<22> ECLK_B<21> ECLK_B<22> WL_O<351> WL_O<350> WL_O<349> WL_O<348> 
+ WL_O<347> WL_O<346> WL_O<345> WL_O<344> WL_O<343> WL_O<342> WL_O<341> 
+ WL_O<340> WL_O<339> WL_O<338> WL_O<337> WL_O<336> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<20> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<20> ECLK_H<20> 
+ ECLK_H<21> ECLK_B<20> ECLK_B<21> WL_O<335> WL_O<334> WL_O<333> WL_O<332> 
+ WL_O<331> WL_O<330> WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> 
+ WL_O<324> WL_O<323> WL_O<322> WL_O<321> WL_O<320> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<19> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<19> ECLK_H<19> 
+ ECLK_H<20> ECLK_B<19> ECLK_B<20> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<18> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<18> ECLK_H<18> 
+ ECLK_H<19> ECLK_B<18> ECLK_B<19> WL_O<303> WL_O<302> WL_O<301> WL_O<300> 
+ WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> WL_O<294> WL_O<293> 
+ WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<17> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<17> ECLK_H<17> 
+ ECLK_H<18> ECLK_B<17> ECLK_B<18> WL_O<287> WL_O<286> WL_O<285> WL_O<284> 
+ WL_O<283> WL_O<282> WL_O<281> WL_O<280> WL_O<279> WL_O<278> WL_O<277> 
+ WL_O<276> WL_O<275> WL_O<274> WL_O<273> WL_O<272> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<16> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<16> ECLK_H<16> 
+ ECLK_H<17> ECLK_B<16> ECLK_B<17> WL_O<271> WL_O<270> WL_O<269> WL_O<268> 
+ WL_O<267> WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> 
+ WL_O<260> WL_O<259> WL_O<258> WL_O<257> WL_O<256> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XDEC10<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<30> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<26> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<22> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<18> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC01<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<29> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<25> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<21> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<17> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XL2<258> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<257> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<256> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<255> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<254> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<253> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<252> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<251> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<250> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<249> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<248> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<247> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<246> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<245> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<244> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<243> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<242> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<241> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<240> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<239> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<238> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<237> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<236> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<235> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<234> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<233> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<232> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<231> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<230> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<229> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<228> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<227> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<226> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<225> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<224> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<223> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<222> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<221> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<220> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<219> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<218> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<217> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<216> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<215> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<214> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<213> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<212> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<211> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<210> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<209> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<208> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<207> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<206> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<205> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<204> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<203> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<202> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<201> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<200> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<199> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<198> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<197> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<196> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<195> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<194> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<193> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<192> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<191> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<190> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<189> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<188> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<187> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<186> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<185> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<184> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<183> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<182> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<181> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<180> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<179> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<178> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<177> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<176> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<175> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<174> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<173> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<172> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<171> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<170> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<169> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<168> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<167> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<166> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<165> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<164> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<163> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<162> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<161> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<160> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<159> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<158> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<157> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<156> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<155> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<154> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<153> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<152> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<151> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<150> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<149> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<148> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<147> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<146> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<145> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<144> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<143> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<142> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<141> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<140> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<139> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<138> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<137> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<136> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<135> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<134> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<133> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC00<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<28> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<24> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<20> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<16> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC11<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<31> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<27> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<23> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<19> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XI0 ADDR_N_I<9> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWREG9 ACLK_N_I ADDR_I<8> ADDR_I<7> ADDR_I<6> ADDR_I<5> 
+ ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<8> ADDR_N_O<7> 
+ ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> 
+ ADDR_N_O<0> BIST_ADDR_I<8> BIST_ADDR_I<7> BIST_ADDR_I<6> BIST_ADDR_I<5> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XDFF<8> BIST_EN_I BIST_ADDR_I<8> ACLK_N_I ADDR_I<8> q_int<8> net04<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net04<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net04<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net04<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net04<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net04<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net04<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net04<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net04<8> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDRV<8> qn_int<8> ADDR_N_O<8> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XINV<8> q_int<8> qn_int<8> VDD VSS / RSC_IHPSG13_CINVX2
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_2P_DLY_MUX A SEL Z VDD VSS
XI11 net4 Z VDD VSS / RSC_IHPSG13_CINVX2
XI8 A D<3> SEL net4 VDD VSS / RSC_IHPSG13_MX2IX1
XI20<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1
XI20<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_CTRL ACLK_N BIST_CK_I BIST_CS_I BIST_EN BIST_RE_I 
+ BIST_WE_I B_TIEL_O CK_I CS_I DCLK ECLK PULSE_H PULSE_L PULSE_O RCLK RE_I 
+ ROW_CS WCLK WE_I VDD VSS
XI17 ck_regs we col_we VDD VSS / RSC_IHPSG13_DFNQX2
XI16 ck_regs re col_re VDD VSS / RSC_IHPSG13_DFNQX2
XI18 ck_regs cs net7 VDD VSS / RSC_IHPSG13_DFNQX2
XI71 ACLK_N net012 PULSE_O VDD VSS / RSC_IHPSG13_DFNQX2
XI77 col_we net017 net016 VDD VSS / RSC_IHPSG13_CNAND2X2
XI76 col_re net017 net018 VDD VSS / RSC_IHPSG13_CNAND2X2
XI15 ck_dly WEorREandCS aclk VDD VSS / RSC_IHPSG13_CGATEPX4
XI14 ck WEandCS DCLK VDD VSS / RSC_IHPSG13_CGATEPX4
XI60 net7 ROW_CS VDD VSS / RSC_IHPSG13_CBUFX8
XI73 PULSE_O net012 VDD VSS / RSC_IHPSG13_CINVX2
XI8 net017 net8 VDD VSS / RSC_IHPSG13_CINVX2
XCAPS4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XCAPS4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XBM_TIEL B_TIEL_O VDD VSS / RSC_IHPSG13_TIEL
XI64 ck ck_dly VDD VSS / RSC_IHPSG13_CDLYX2
XI86 CS_I BIST_CS_I BIST_EN cs VDD VSS / RSC_IHPSG13_MX2X2
XI87 CK_I BIST_CK_I BIST_EN ck VDD VSS / RSC_IHPSG13_MX2X2
XI85 WE_I BIST_WE_I BIST_EN we VDD VSS / RSC_IHPSG13_MX2X2
XI84 RE_I BIST_RE_I BIST_EN re VDD VSS / RSC_IHPSG13_MX2X2
XI48 ck_dly ck_regs VDD VSS / RSC_IHPSG13_CINVX4
XI81 net016 WCLK VDD VSS / RSC_IHPSG13_CINVX4
XI80 net018 RCLK VDD VSS / RSC_IHPSG13_CINVX4
XI78 net8 net020 VDD VSS / RSC_IHPSG13_CINVX4
XCAPS8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XCAPS8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI6 PULSE_L PULSE_H net017 VDD VSS / RSC_IHPSG13_XOR2X2
XI22 we cs WEandCS VDD VSS / RSC_IHPSG13_AND2X2
XI79 net020 ECLK VDD VSS / RSC_IHPSG13_CINVX8
XI63 aclk ACLK_N VDD VSS / RSC_IHPSG13_CINVX8
XI21 re we cs WEorREandCS VDD VSS / RSC_IHPSG13_OA12X1
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDEC5 ACLK_N ADDR<4> ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<4> BIST_ADDR<3> 
+ BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<4> BIST_EN_I BIST_ADDR<4> ACLK_N ADDR<4> addr_int<1> net13<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int<0> net13<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net13<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net13<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net13<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI15<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI15<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> addr_int<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_CBUFX2
XI13<0> addr_int<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XI14<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI14<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_BLDRV A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> 
+ A_SEL_P<1> A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> 
+ B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> 
+ B_SEL_P<2> B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS
MA_CWN<3> A_BLC<3> A_BLC_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<2> A_BLC<2> A_BLC_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<1> A_BLC<1> A_BLC_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CWN<0> A_BLC<0> A_BLC_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<3> A_BLT<3> A_BLT_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<2> A_BLT<2> A_BLT_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<1> A_BLT<1> A_BLT_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_TWN<0> A_BLT<0> A_BLT_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<3> B_BLT<3> B_BLT_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<2> B_BLT<2> B_BLT_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<1> B_BLT<1> B_BLT_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_TWN<0> B_BLT<0> B_BLT_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<3> B_BLC<3> B_BLC_NMOS_DRIVE<3> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<2> B_BLC<2> B_BLC_NMOS_DRIVE<2> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<1> B_BLC<1> B_BLC_NMOS_DRIVE<1> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MB_CWN<0> B_BLC<0> B_BLC_NMOS_DRIVE<0> VSS VSS nmos m=1 
+ w=4.82u l=130.00n ng=2 nrd=0 nrs=0
MA_CPR<3> A_BLC<3> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<2> A_BLC<2> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<1> A_BLC<1> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_CPR<0> A_BLC<0> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TWP<3> A_BLT<3> A_BLT_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<2> A_BLT<2> A_BLT_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<1> A_BLT<1> A_BLT_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TWP<0> A_BLT<0> A_BLT_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<3> A_BLC<3> A_BLC_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<2> A_BLC<2> A_BLC_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<1> A_BLC<1> A_BLC_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CWP<0> A_BLC<0> A_BLC_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TPR<3> A_BLT<3> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<2> A_BLT<2> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<1> A_BLT<1> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TPR<0> A_BLT<0> A_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MA_TSP<3> A_BLT_SEL A_SEL_N<3> A_BLT<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<2> A_BLT_SEL A_SEL_N<2> A_BLT<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<1> A_BLT_SEL A_SEL_N<1> A_BLT<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_TSP<0> A_BLT_SEL A_SEL_N<0> A_BLT<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<3> A_BLC_SEL A_SEL_N<3> A_BLC<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<2> A_BLC_SEL A_SEL_N<2> A_BLC<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<1> A_BLC_SEL A_SEL_N<1> A_BLC<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MA_CSP<0> A_BLC_SEL A_SEL_N<0> A_BLC<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<3> B_BLC<3> B_BLC_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<2> B_BLC<2> B_BLC_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<1> B_BLC<1> B_BLC_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CWP<0> B_BLC<0> B_BLC_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<3> B_BLT<3> B_BLT_PMOS_DRIVE<3> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<2> B_BLT<2> B_BLT_PMOS_DRIVE<2> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<1> B_BLT<1> B_BLT_PMOS_DRIVE<1> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TWP<0> B_BLT<0> B_BLT_PMOS_DRIVE<0> VDD VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<3> B_BLT_SEL B_SEL_N<3> B_BLT<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<2> B_BLT_SEL B_SEL_N<2> B_BLT<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<1> B_BLT_SEL B_SEL_N<1> B_BLT<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TSP<0> B_BLT_SEL B_SEL_N<0> B_BLT<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_TPR<3> B_BLT<3> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<2> B_BLT<2> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<1> B_BLT<1> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_TPR<0> B_BLT<0> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CSP<3> B_BLC_SEL B_SEL_N<3> B_BLC<3> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<2> B_BLC_SEL B_SEL_N<2> B_BLC<2> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<1> B_BLC_SEL B_SEL_N<1> B_BLC<1> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CSP<0> B_BLC_SEL B_SEL_N<0> B_BLC<0> VDD pmos m=1 w=1.5u 
+ l=130.00n ng=1 nrd=0 nrs=0
MB_CPR<3> B_BLC<3> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<2> B_BLC<2> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<1> B_BLC<1> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
MB_CPR<0> B_BLC<0> B_PRE_N VDD VDD pmos m=1 w=3.000u l=130.00n 
+ ng=2 nrd=0 nrs=0
XA_SEL<3> A_SEL_P<3> A_SEL_N<3> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<2> A_SEL_P<2> A_SEL_N<2> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<1> A_SEL_P<1> A_SEL_N<1> VDD VSS / RSC_IHPSG13_INVX2
XA_SEL<0> A_SEL_P<0> A_SEL_N<0> VDD VSS / RSC_IHPSG13_INVX2
XA_CINV<3> A_BLT_PMOS_DRIVE<3> A_BLC_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<2> A_BLT_PMOS_DRIVE<2> A_BLC_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<1> A_BLT_PMOS_DRIVE<1> A_BLC_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_CINV<0> A_BLT_PMOS_DRIVE<0> A_BLC_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<3> A_BLC_PMOS_DRIVE<3> A_BLT_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<2> A_BLC_PMOS_DRIVE<2> A_BLT_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<1> A_BLC_PMOS_DRIVE<1> A_BLT_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TINV<0> A_BLC_PMOS_DRIVE<0> A_BLT_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_SEL<3> B_SEL_P<3> B_SEL_N<3> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<2> B_SEL_P<2> B_SEL_N<2> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<1> B_SEL_P<1> B_SEL_N<1> VDD VSS / RSC_IHPSG13_INVX2
XB_SEL<0> B_SEL_P<0> B_SEL_N<0> VDD VSS / RSC_IHPSG13_INVX2
XB_TINV<3> B_BLC_PMOS_DRIVE<3> B_BLT_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<2> B_BLC_PMOS_DRIVE<2> B_BLT_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<1> B_BLC_PMOS_DRIVE<1> B_BLT_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_TINV<0> B_BLC_PMOS_DRIVE<0> B_BLT_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<3> B_BLT_PMOS_DRIVE<3> B_BLC_NMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<2> B_BLT_PMOS_DRIVE<2> B_BLC_NMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<1> B_BLT_PMOS_DRIVE<1> B_BLC_NMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_INVX2
XB_CINV<0> B_BLT_PMOS_DRIVE<0> B_BLC_NMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_INVX2
XA_TDEC<3> A_SEL_P<3> A_WR_ONE A_BLT_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<2> A_SEL_P<2> A_WR_ONE A_BLT_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<1> A_SEL_P<1> A_WR_ONE A_BLT_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_TDEC<0> A_SEL_P<0> A_WR_ONE A_BLT_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<3> A_SEL_P<3> A_WR_ZERO A_BLC_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<2> A_SEL_P<2> A_WR_ZERO A_BLC_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<1> A_SEL_P<1> A_WR_ZERO A_BLC_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XA_CDEC<0> A_SEL_P<0> A_WR_ZERO A_BLC_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<3> B_SEL_P<3> B_WR_ZERO B_BLC_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<2> B_SEL_P<2> B_WR_ZERO B_BLC_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<1> B_SEL_P<1> B_WR_ZERO B_BLC_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_CDEC<0> B_SEL_P<0> B_WR_ZERO B_BLC_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<3> B_SEL_P<3> B_WR_ONE B_BLT_PMOS_DRIVE<3> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<2> B_SEL_P<2> B_WR_ONE B_BLT_PMOS_DRIVE<2> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<1> B_SEL_P<1> B_WR_ONE B_BLT_PMOS_DRIVE<1> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
XB_TDEC<0> B_SEL_P<0> B_WR_ONE B_BLT_PMOS_DRIVE<0> VDD VSS / 
+ RSC_IHPSG13_NAND2X2
.ENDS
.SUBCKT RSC_IHPSG13_AND2X6 A B Z VDD VSS
MN3 Z net6 VSS VSS nmos m=1 w=2.94u l=130.00n ng=3 nrd=0 nrs=0
MN4 net9 B VSS VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MN6 net6 A net9 VSS nmos m=1 w=500.0n l=130.00n ng=1 nrd=0 nrs=0
MP2 Z net6 VDD VDD pmos m=1 w=4.86u l=130.00n ng=3 nrd=0 nrs=0
MP0 net6 B VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
MP1 net6 A VDD VDD pmos m=1 w=860.00n l=130.00n ng=1 nrd=0 
+ nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLCTRL5 A_ADDR_COL<1> A_ADDR_COL<0> A_ADDR_DEC<7> 
+ A_ADDR_DEC<6> A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<31> 
+ A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> 
+ A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> 
+ A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> 
+ A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> 
+ A_BLC<1> A_BLC<0> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> 
+ A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> 
+ A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> 
+ A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_COL<1> B_ADDR_COL<0> 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> 
+ B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I 
+ B_BIST_EN_I B_BLC<31> B_BLC<30> B_BLC<29> B_BLC<28> B_BLC<27> B_BLC<26> 
+ B_BLC<25> B_BLC<24> B_BLC<23> B_BLC<22> B_BLC<21> B_BLC<20> B_BLC<19> 
+ B_BLC<18> B_BLC<17> B_BLC<16> B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> 
+ B_BLC<11> B_BLC<10> B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> 
+ B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<31> B_BLT<30> B_BLT<29> B_BLT<28> 
+ B_BLT<27> B_BLT<26> B_BLT<25> B_BLT<24> B_BLT<23> B_BLT<22> B_BLT<21> 
+ B_BLT<20> B_BLT<19> B_BLT<18> B_BLT<17> B_BLT<16> B_BLT<15> B_BLT<14> 
+ B_BLT<13> B_BLT<12> B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> 
+ B_BLT<5> B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L 
+ B_DCLK_B_R B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L 
+ B_RCLK_R B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_I80<1> B_WCLK_B_L B_RCLK_B_L B_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XB_I80<0> B_WCLK_B_L B_RCLK_B_L B_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<1> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<0> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XI_FILL4<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XB_INV<6> B_N1<1> B_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<5> B_N0<1> B_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<4> B_N0<0> B_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<3> B_ADDR_COL<1> B_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<2> B_ADDR_COL<1> B_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<1> B_ADDR_COL<0> B_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<0> B_ADDR_COL<0> B_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<6> A_N1<1> A_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<5> A_N0<1> A_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<4> A_N0<0> A_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<3> A_ADDR_COL<1> A_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<2> A_ADDR_COL<1> A_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_ADDR_COL<0> A_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL<0> A_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XB_I81<3> B_W_nor_R<1> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<2> B_W_nor_R<1> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<1> B_W_nor_R<0> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<0> B_W_nor_R<0> B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<3> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<2> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XI_FILL8<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XAB_BLMUX<7> A_BLC<31> A_BLC<30> A_BLC<29> A_BLC<28> A_BLC_SEL A_BLT<31> 
+ A_BLT<30> A_BLT<29> A_BLT<28> A_BLT_SEL A_PRE_N A_SEL_P<31> A_SEL_P<30> 
+ A_SEL_P<29> A_SEL_P<28> A_WR_ONE A_WR_ZERO B_BLC<31> B_BLC<30> B_BLC<29> 
+ B_BLC<28> B_BLC_SEL B_BLT<31> B_BLT<30> B_BLT<29> B_BLT<28> B_BLT_SEL 
+ B_PRE_N B_SEL_P<31> B_SEL_P<30> B_SEL_P<29> B_SEL_P<28> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<6> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> A_BLC_SEL A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT_SEL A_PRE_N A_SEL_P<27> A_SEL_P<26> 
+ A_SEL_P<25> A_SEL_P<24> A_WR_ONE A_WR_ZERO B_BLC<27> B_BLC<26> B_BLC<25> 
+ B_BLC<24> B_BLC_SEL B_BLT<27> B_BLT<26> B_BLT<25> B_BLT<24> B_BLT_SEL 
+ B_PRE_N B_SEL_P<27> B_SEL_P<26> B_SEL_P<25> B_SEL_P<24> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<5> A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC_SEL A_BLT<23> 
+ A_BLT<22> A_BLT<21> A_BLT<20> A_BLT_SEL A_PRE_N A_SEL_P<23> A_SEL_P<22> 
+ A_SEL_P<21> A_SEL_P<20> A_WR_ONE A_WR_ZERO B_BLC<23> B_BLC<22> B_BLC<21> 
+ B_BLC<20> B_BLC_SEL B_BLT<23> B_BLT<22> B_BLT<21> B_BLT<20> B_BLT_SEL 
+ B_PRE_N B_SEL_P<23> B_SEL_P<22> B_SEL_P<21> B_SEL_P<20> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<4> A_BLC<19> A_BLC<18> A_BLC<17> A_BLC<16> A_BLC_SEL A_BLT<19> 
+ A_BLT<18> A_BLT<17> A_BLT<16> A_BLT_SEL A_PRE_N A_SEL_P<19> A_SEL_P<18> 
+ A_SEL_P<17> A_SEL_P<16> A_WR_ONE A_WR_ZERO B_BLC<19> B_BLC<18> B_BLC<17> 
+ B_BLC<16> B_BLC_SEL B_BLT<19> B_BLT<18> B_BLT<17> B_BLT<16> B_BLT_SEL 
+ B_PRE_N B_SEL_P<19> B_SEL_P<18> B_SEL_P<17> B_SEL_P<16> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<3> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC_SEL A_BLT<15> 
+ A_BLT<14> A_BLT<13> A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<15> A_SEL_P<14> 
+ A_SEL_P<13> A_SEL_P<12> A_WR_ONE A_WR_ZERO B_BLC<15> B_BLC<14> B_BLC<13> 
+ B_BLC<12> B_BLC_SEL B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT_SEL 
+ B_PRE_N B_SEL_P<15> B_SEL_P<14> B_SEL_P<13> B_SEL_P<12> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<2> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC_SEL A_BLT<11> 
+ A_BLT<10> A_BLT<9> A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<11> A_SEL_P<10> 
+ A_SEL_P<9> A_SEL_P<8> A_WR_ONE A_WR_ZERO B_BLC<11> B_BLC<10> B_BLC<9> 
+ B_BLC<8> B_BLC_SEL B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT_SEL B_PRE_N 
+ B_SEL_P<11> B_SEL_P<10> B_SEL_P<9> B_SEL_P<8> B_WR_ONE B_WR_ZERO VDD 
+ VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<7> A_SEL_P<6> A_SEL_P<5> 
+ A_SEL_P<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC_SEL 
+ B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N B_SEL_P<7> B_SEL_P<6> 
+ B_SEL_P<5> B_SEL_P<4> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> A_SEL_P<1> 
+ A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLC_SEL 
+ B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> B_SEL_P<2> 
+ B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BLDRV
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<31> net041<0> B_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<30> net041<1> B_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<29> net041<2> B_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<28> net041<3> B_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<27> net041<4> B_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<26> net041<5> B_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<25> net041<6> B_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<24> net041<7> B_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<23> net041<8> B_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<22> net041<9> B_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<21> net041<10> B_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<20> net041<11> B_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<19> net041<12> B_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<18> net041<13> B_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<17> net041<14> B_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<16> net041<15> B_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<15> net041<16> B_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<14> net041<17> B_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<13> net041<18> B_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<12> net041<19> B_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<11> net041<20> B_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<10> net041<21> B_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<9> net041<22> B_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<8> net041<23> B_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<7> net041<24> B_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<6> net041<25> B_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<5> net041<26> B_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<4> net041<27> B_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<3> net041<28> B_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<2> net041<29> B_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<1> net041<30> B_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<0> net041<31> B_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<31> net23<0> A_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<30> net23<1> A_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<29> net23<2> A_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<28> net23<3> A_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<27> net23<4> A_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<26> net23<5> A_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<25> net23<6> A_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<24> net23<7> A_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<23> net23<8> A_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<22> net23<9> A_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<21> net23<10> A_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<20> net23<11> A_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<19> net23<12> A_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<18> net23<13> A_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<17> net23<14> A_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<16> net23<15> A_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<15> net23<16> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<17> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<18> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<19> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<20> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<21> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<22> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<23> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<24> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<25> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<26> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<27> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<28> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<29> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<30> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<31> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net042 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net043 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net21 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_DEC3<31> B_P1<1> B_P0<1> B_ADDR_DEC<7> net041<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<30> B_P1<1> B_P0<1> B_ADDR_DEC<6> net041<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<29> B_P1<1> B_P0<1> B_ADDR_DEC<5> net041<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<28> B_P1<1> B_P0<1> B_ADDR_DEC<4> net041<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<27> B_P1<1> B_P0<1> B_ADDR_DEC<3> net041<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<26> B_P1<1> B_P0<1> B_ADDR_DEC<2> net041<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<25> B_P1<1> B_P0<1> B_ADDR_DEC<1> net041<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<24> B_P1<1> B_P0<1> B_ADDR_DEC<0> net041<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<23> B_P1<1> B_N0<1> B_ADDR_DEC<7> net041<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<22> B_P1<1> B_N0<1> B_ADDR_DEC<6> net041<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<21> B_P1<1> B_N0<1> B_ADDR_DEC<5> net041<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<20> B_P1<1> B_N0<1> B_ADDR_DEC<4> net041<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<19> B_P1<1> B_N0<1> B_ADDR_DEC<3> net041<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<18> B_P1<1> B_N0<1> B_ADDR_DEC<2> net041<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<17> B_P1<1> B_N0<1> B_ADDR_DEC<1> net041<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<16> B_P1<1> B_N0<1> B_ADDR_DEC<0> net041<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<15> B_N1<0> B_P0<0> B_ADDR_DEC<7> net041<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<14> B_N1<0> B_P0<0> B_ADDR_DEC<6> net041<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<13> B_N1<0> B_P0<0> B_ADDR_DEC<5> net041<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<12> B_N1<0> B_P0<0> B_ADDR_DEC<4> net041<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<11> B_N1<0> B_P0<0> B_ADDR_DEC<3> net041<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<10> B_N1<0> B_P0<0> B_ADDR_DEC<2> net041<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<9> B_N1<0> B_P0<0> B_ADDR_DEC<1> net041<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<8> B_N1<0> B_P0<0> B_ADDR_DEC<0> net041<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<7> B_N1<0> B_N0<0> B_ADDR_DEC<7> net041<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<6> B_N1<0> B_N0<0> B_ADDR_DEC<6> net041<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<5> B_N1<0> B_N0<0> B_ADDR_DEC<5> net041<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<4> B_N1<0> B_N0<0> B_ADDR_DEC<4> net041<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<3> B_N1<0> B_N0<0> B_ADDR_DEC<3> net041<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<2> B_N1<0> B_N0<0> B_ADDR_DEC<2> net041<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<1> B_N1<0> B_N0<0> B_ADDR_DEC<1> net041<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_DEC3<0> B_N1<0> B_N0<0> B_ADDR_DEC<0> net041<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<31> A_P1<1> A_P0<1> A_ADDR_DEC<7> net23<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<30> A_P1<1> A_P0<1> A_ADDR_DEC<6> net23<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<29> A_P1<1> A_P0<1> A_ADDR_DEC<5> net23<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<28> A_P1<1> A_P0<1> A_ADDR_DEC<4> net23<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<27> A_P1<1> A_P0<1> A_ADDR_DEC<3> net23<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<26> A_P1<1> A_P0<1> A_ADDR_DEC<2> net23<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<25> A_P1<1> A_P0<1> A_ADDR_DEC<1> net23<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<24> A_P1<1> A_P0<1> A_ADDR_DEC<0> net23<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<23> A_P1<1> A_N0<1> A_ADDR_DEC<7> net23<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<22> A_P1<1> A_N0<1> A_ADDR_DEC<6> net23<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<21> A_P1<1> A_N0<1> A_ADDR_DEC<5> net23<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<20> A_P1<1> A_N0<1> A_ADDR_DEC<4> net23<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<19> A_P1<1> A_N0<1> A_ADDR_DEC<3> net23<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<18> A_P1<1> A_N0<1> A_ADDR_DEC<2> net23<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<17> A_P1<1> A_N0<1> A_ADDR_DEC<1> net23<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<16> A_P1<1> A_N0<1> A_ADDR_DEC<0> net23<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<15> A_N1<0> A_P0<0> A_ADDR_DEC<7> net23<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<14> A_N1<0> A_P0<0> A_ADDR_DEC<6> net23<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<13> A_N1<0> A_P0<0> A_ADDR_DEC<5> net23<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<12> A_N1<0> A_P0<0> A_ADDR_DEC<4> net23<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<11> A_N1<0> A_P0<0> A_ADDR_DEC<3> net23<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<10> A_N1<0> A_P0<0> A_ADDR_DEC<2> net23<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<9> A_N1<0> A_P0<0> A_ADDR_DEC<1> net23<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<8> A_N1<0> A_P0<0> A_ADDR_DEC<0> net23<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<7> A_N1<0> A_N0<0> A_ADDR_DEC<7> net23<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<6> A_N1<0> A_N0<0> A_ADDR_DEC<6> net23<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<5> A_N1<0> A_N0<0> A_ADDR_DEC<5> net23<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<4> A_N1<0> A_N0<0> A_ADDR_DEC<4> net23<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<3> A_N1<0> A_N0<0> A_ADDR_DEC<3> net23<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<2> A_N1<0> A_N0<0> A_ADDR_DEC<2> net23<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<1> A_N1<0> A_N0<0> A_ADDR_DEC<1> net23<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<0> A_N1<0> A_N0<0> A_ADDR_DEC<0> net23<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDRV13_FILL4 VDD VSS
XI0<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RSC_IHPSG13_CBUFX16 A Z VDD VSS
MN0 net4 A VSS VSS nmos m=1 w=2.115u l=130.00n ng=3 nrd=0 nrs=0
MN1 Z net4 VSS VSS nmos m=1 w=5.64u l=130.00n ng=8 nrd=0 nrs=0
MP1 Z net4 VDD VDD pmos m=1 w=13.000u l=130.00n ng=8 nrd=0 
+ nrs=0
MP0 net4 A VDD VDD pmos m=1 w=4.89u l=130.00n ng=3 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDRV13X16 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX16 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=12.96u l=130.00n ng=8 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_WLDRV16X16 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX16
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDRV13X4 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1 VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_WLDRV16X4 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX4
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWDEC8 ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> 
+ ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<255> 
+ WL_O<254> WL_O<253> WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> 
+ WL_O<247> WL_O<246> WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> 
+ WL_O<240> WL_O<239> WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> 
+ WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> 
+ WL_O<226> WL_O<225> WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> 
+ WL_O<205> WL_O<204> WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> 
+ WL_O<198> WL_O<197> WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> 
+ WL_O<191> WL_O<190> WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> 
+ WL_O<184> WL_O<183> WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> 
+ WL_O<177> WL_O<176> WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> 
+ WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> 
+ WL_O<163> WL_O<162> WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> 
+ WL_O<156> WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> 
+ WL_O<149> WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> 
+ WL_O<142> WL_O<141> WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> 
+ WL_O<135> WL_O<134> WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> 
+ WL_O<128> WL_O<127> WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> 
+ WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> 
+ WL_O<114> WL_O<113> WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> 
+ WL_O<92> WL_O<91> WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> 
+ WL_O<84> WL_O<83> WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> 
+ WL_O<76> WL_O<75> WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> 
+ WL_O<68> WL_O<67> WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> 
+ WL_O<60> WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> 
+ WL_O<52> WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> 
+ WL_O<44> WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> 
+ WL_O<36> WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> 
+ WL_O<28> WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> 
+ WL_O<20> WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> 
+ WL_O<12> WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> 
+ WL_O<3> WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XDEC10<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC00<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC01<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWREG8 ACLK_N_I ADDR_I<7> ADDR_I<6> ADDR_I<5> ADDR_I<4> 
+ ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<7> ADDR_N_O<6> ADDR_N_O<5> 
+ ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<7> 
+ BIST_ADDR_I<6> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> 
+ BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI10 VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDEC4 ACLK_N ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<3> BIST_ADDR<2> 
+ BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int net12<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net12<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net12<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net12<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI14 addr_int ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI15 ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLCTRL4 A_ADDR_COL A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<15> A_BLC<14> 
+ A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> 
+ A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<15> A_BLT<14> 
+ A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L 
+ A_DCLK_B_R A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L 
+ A_RCLK_R A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_COL 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> 
+ B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I 
+ B_BIST_EN_I B_BLC<15> B_BLC<14> B_BLC<13> B_BLC<12> B_BLC<11> B_BLC<10> 
+ B_BLC<9> B_BLC<8> B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC<3> B_BLC<2> 
+ B_BLC<1> B_BLC<0> B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT<11> 
+ B_BLT<10> B_BLT<9> B_BLT<8> B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT<3> 
+ B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L B_DCLK_B_R B_DCLK_L B_DCLK_R 
+ B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L B_RCLK_R B_TIEH_O B_WCLK_B_L 
+ B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_I80 B_RCLK_B_L B_WCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_RCLK_B_L A_WCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X4
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X4
XI_FILL4<26> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<25> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<24> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<23> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<22> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<21> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<20> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<19> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<18> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<17> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<1> B_N0 B_P0 VDD VSS / RSC_IHPSG13_CINVX4
XB_INV<0> B_ADDR_COL B_N0 VDD VSS / RSC_IHPSG13_CINVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_N0 A_P0 VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL A_N0 VDD VSS / RSC_IHPSG13_CINVX4
XB_I81<1> net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_I81<0> net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XAB_BLMUX<3> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC_SEL A_BLT<15> 
+ A_BLT<14> A_BLT<13> A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<15> A_SEL_P<14> 
+ A_SEL_P<13> A_SEL_P<12> A_WR_ONE A_WR_ZERO B_BLC<15> B_BLC<14> B_BLC<13> 
+ B_BLC<12> B_BLC_SEL B_BLT<15> B_BLT<14> B_BLT<13> B_BLT<12> B_BLT_SEL 
+ B_PRE_N B_SEL_P<15> B_SEL_P<14> B_SEL_P<13> B_SEL_P<12> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<2> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC_SEL A_BLT<11> 
+ A_BLT<10> A_BLT<9> A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<11> A_SEL_P<10> 
+ A_SEL_P<9> A_SEL_P<8> A_WR_ONE A_WR_ZERO B_BLC<11> B_BLC<10> B_BLC<9> 
+ B_BLC<8> B_BLC_SEL B_BLT<11> B_BLT<10> B_BLT<9> B_BLT<8> B_BLT_SEL B_PRE_N 
+ B_SEL_P<11> B_SEL_P<10> B_SEL_P<9> B_SEL_P<8> B_WR_ONE B_WR_ZERO VDD 
+ VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<7> A_SEL_P<6> A_SEL_P<5> 
+ A_SEL_P<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> B_BLC<4> B_BLC_SEL 
+ B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N B_SEL_P<7> B_SEL_P<6> 
+ B_SEL_P<5> B_SEL_P<4> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<3> A_SEL_P<2> A_SEL_P<1> 
+ A_SEL_P<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLC_SEL 
+ B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N B_SEL_P<3> B_SEL_P<2> 
+ B_SEL_P<1> B_SEL_P<0> B_WR_ONE B_WR_ZERO VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_BLDRV
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net046 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net045 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net24 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3INV<15> net23<0> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<1> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<2> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<3> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<4> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<5> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<6> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<7> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<8> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<9> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<10> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<11> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<12> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<13> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<14> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<15> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<15> net044<0> B_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<14> net044<1> B_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<13> net044<2> B_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<12> net044<3> B_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<11> net044<4> B_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<10> net044<5> B_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<9> net044<6> B_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<8> net044<7> B_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<7> net044<8> B_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<6> net044<9> B_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<5> net044<10> B_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<4> net044<11> B_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<3> net044<12> B_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<2> net044<13> B_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<1> net044<14> B_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XB_DEC3INV<0> net044<15> B_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XI_FILL8<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_DEC3<15> A_P0 A_ADDR_DEC<7> net23<0> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<14> A_P0 A_ADDR_DEC<6> net23<1> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<13> A_P0 A_ADDR_DEC<5> net23<2> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<12> A_P0 A_ADDR_DEC<4> net23<3> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<11> A_P0 A_ADDR_DEC<3> net23<4> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<10> A_P0 A_ADDR_DEC<2> net23<5> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<9> A_P0 A_ADDR_DEC<1> net23<6> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<8> A_P0 A_ADDR_DEC<0> net23<7> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<7> A_N0 A_ADDR_DEC<7> net23<8> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<6> A_N0 A_ADDR_DEC<6> net23<9> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<5> A_N0 A_ADDR_DEC<5> net23<10> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<4> A_N0 A_ADDR_DEC<4> net23<11> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<3> A_N0 A_ADDR_DEC<3> net23<12> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<2> A_N0 A_ADDR_DEC<2> net23<13> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<1> A_N0 A_ADDR_DEC<1> net23<14> VDD VSS / RSC_IHPSG13_NAND2X2
XA_DEC3<0> A_N0 A_ADDR_DEC<0> net23<15> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<15> B_P0 B_ADDR_DEC<7> net044<0> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<14> B_P0 B_ADDR_DEC<6> net044<1> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<13> B_P0 B_ADDR_DEC<5> net044<2> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<12> B_P0 B_ADDR_DEC<4> net044<3> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<11> B_P0 B_ADDR_DEC<3> net044<4> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<10> B_P0 B_ADDR_DEC<2> net044<5> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<9> B_P0 B_ADDR_DEC<1> net044<6> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<8> B_P0 B_ADDR_DEC<0> net044<7> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<7> B_N0 B_ADDR_DEC<7> net044<8> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<6> B_N0 B_ADDR_DEC<6> net044<9> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<5> B_N0 B_ADDR_DEC<5> net044<10> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<4> B_N0 B_ADDR_DEC<4> net044<11> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<3> B_N0 B_ADDR_DEC<3> net044<12> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<2> B_N0 B_ADDR_DEC<2> net044<13> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<1> B_N0 B_ADDR_DEC<1> net044<14> VDD VSS / RSC_IHPSG13_NAND2X2
XB_DEC3<0> B_N0 B_ADDR_DEC<0> net044<15> VDD VSS / RSC_IHPSG13_NAND2X2
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWDEC5 ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> 
+ ADDR_N_I<0> CS_I ECLK_I WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0 ADDR_N_I<5> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWREG5 ACLK_N_I ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> 
+ ADDR_I<0> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDEC3 ACLK_N ADDR<2> ADDR<1> ADDR<0> ADDR_COL<1> 
+ ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> 
+ ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> 
+ BIST_EN_I VDD VSS
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net13<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net13<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net13<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI15<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI15<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI13<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XI17<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_DFPQD_MSAFFX2P CP DN DP QN QP VDD VSS
XI_AMP CP DN DP QN QP VDD VSS / RSC_IHPSG13_DFPQD_MSAFFX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLCTRL3 A_ADDR_DEC<7> A_ADDR_DEC<6> A_ADDR_DEC<5> 
+ A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> A_ADDR_DEC<0> 
+ A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> 
+ A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> 
+ A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R A_DCLK_L 
+ A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R A_TIEH_O 
+ A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_DEC<7> B_ADDR_DEC<6> 
+ B_ADDR_DEC<5> B_ADDR_DEC<4> B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> 
+ B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I B_BIST_EN_I B_BLC<7> B_BLC<6> B_BLC<5> 
+ B_BLC<4> B_BLC<3> B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<7> B_BLT<6> B_BLT<5> 
+ B_BLT<4> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I B_DCLK_B_L B_DCLK_B_R 
+ B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R B_RCLK_L B_RCLK_R 
+ B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD VSS
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net044 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net043 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XI_FILL8<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI_FILL8<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XB_I51 net037 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XB_I44 B_BM_N B_WCLK_B_L B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net037 net038 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2P
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2P
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XAB_BLMUX<1> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC_SEL A_BLT<7> A_BLT<6> 
+ A_BLT<5> A_BLT<4> A_BLT_SEL A_PRE_N A_ADDR_DEC<7> A_ADDR_DEC<6> 
+ A_ADDR_DEC<5> A_ADDR_DEC<4> A_WR_ONE A_WR_ZERO B_BLC<7> B_BLC<6> B_BLC<5> 
+ B_BLC<4> B_BLC_SEL B_BLT<7> B_BLT<6> B_BLT<5> B_BLT<4> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<7> B_ADDR_DEC<6> B_ADDR_DEC<5> B_ADDR_DEC<4> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XAB_BLMUX<0> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> 
+ B_BLC<0> B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I80 B_WCLK_B_L B_RCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DO_WRITE_P B_DI_N B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XB_I75 B_DO_WRITE_P B_DI_R B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_WCLK_B_L A_RCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XB_I81 net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XI_FILL4<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI_FILL4<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWDEC6 ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> 
+ ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<63> WL_O<62> WL_O<61> WL_O<60> 
+ WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> 
+ WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> 
+ WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> 
+ WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> 
+ WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> 
+ WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> 
+ WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> 
+ WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC10 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XDEC11 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWREG6 ACLK_N_I ADDR_I<5> ADDR_I<4> ADDR_I<3> ADDR_I<2> 
+ ADDR_I<1> ADDR_I<0> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> 
+ ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDRV13X16 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX16
XI1<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_WLDRV16X16 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX16
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX16
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_DEC01 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC NADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XI2 VDD VSS / RSC_IHPSG13_FILLCAP4
XADDRINV ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_DEC00 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC NADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XADDRINV<1> ADDR<1> NADDR<1> VDD VSS / RSC_IHPSG13_INVX2
XADDRINV<0> ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
XI1 VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWDEC5 ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> 
+ ADDR_N_I<0> CS_I ECLK_I WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XI0 ADDR_N_I<5> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWREG5 ACLK_N_I ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> 
+ ADDR_I<0> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDEC5 ACLK_N ADDR<4> ADDR<3> ADDR<2> ADDR<1> ADDR<0> 
+ ADDR_COL<1> ADDR_COL<0> ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> 
+ ADDR_DEC<3> ADDR_DEC<2> ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<4> BIST_ADDR<3> 
+ BIST_ADDR<2> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI17<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI17<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI13<1> addr_int<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_CBUFX2
XI13<0> addr_int<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_CBUFX2
XDFF<4> BIST_EN_I BIST_ADDR<4> ACLK_N ADDR<4> addr_int<1> net7<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR<3> ACLK_N ADDR<3> addr_int<0> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR<2> ACLK_N ADDR<2> padr_int<2> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net7<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI1<7> PADR<0> PADR<1> PADR<2> addr_n<7> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<6> NADR<0> PADR<1> PADR<2> addr_n<6> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<5> PADR<0> NADR<1> PADR<2> addr_n<5> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<4> NADR<0> NADR<1> PADR<2> addr_n<4> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<3> PADR<0> PADR<1> NADR<2> addr_n<3> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<2> NADR<0> PADR<1> NADR<2> addr_n<2> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<1> PADR<0> NADR<1> NADR<2> addr_n<1> VDD VSS / RSC_IHPSG13_NAND3X2
XI1<0> NADR<0> NADR<1> NADR<2> addr_n<0> VDD VSS / RSC_IHPSG13_NAND3X2
XI15<2> NADR<2> PADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI15<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI15<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<2> padr_int<2> NADR<2> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<7> addr_n<7> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_INVX2
XI2<6> addr_n<6> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_INVX2
XI2<5> addr_n<5> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_INVX2
XI2<4> addr_n<4> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLCTRL5 A_ADDR_COL<1> A_ADDR_COL<0> A_ADDR_DEC<7> 
+ A_ADDR_DEC<6> A_ADDR_DEC<5> A_ADDR_DEC<4> A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<31> 
+ A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> 
+ A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> 
+ A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> 
+ A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> 
+ A_BLC<1> A_BLC<0> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> 
+ A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> 
+ A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> 
+ A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> 
+ A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R VDD VSS
XA_I80<1> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<1> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I80<0> A_WCLK_B_L A_RCLK_B_L A_W_nor_R<0> VDD VSS / 
+ RSC_IHPSG13_AND2X2
XA_I44 A_BM_N A_WCLK_B_L A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XI80<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI80<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_I74<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XA_INV<6> A_N1<1> A_P1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<5> A_N0<1> A_P0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<4> A_N0<0> A_P0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<3> A_ADDR_COL<1> A_N1<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<2> A_ADDR_COL<1> A_N1<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<1> A_ADDR_COL<0> A_N0<1> VDD VSS / RSC_IHPSG13_CINVX4
XA_INV<0> A_ADDR_COL<0> A_N0<0> VDD VSS / RSC_IHPSG13_CINVX4
XA_I81<3> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<2> A_W_nor_R<1> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<1> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81<0> A_W_nor_R<0> A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_BLTMUX<31> A_BLC<31> A_BLC_SEL A_BLT<31> A_BLT_SEL A_PRE_N A_SEL_P<31> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<30> A_BLC<30> A_BLC_SEL A_BLT<30> A_BLT_SEL A_PRE_N A_SEL_P<30> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<29> A_BLC<29> A_BLC_SEL A_BLT<29> A_BLT_SEL A_PRE_N A_SEL_P<29> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<28> A_BLC<28> A_BLC_SEL A_BLT<28> A_BLT_SEL A_PRE_N A_SEL_P<28> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<27> A_BLC<27> A_BLC_SEL A_BLT<27> A_BLT_SEL A_PRE_N A_SEL_P<27> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<26> A_BLC<26> A_BLC_SEL A_BLT<26> A_BLT_SEL A_PRE_N A_SEL_P<26> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<25> A_BLC<25> A_BLC_SEL A_BLT<25> A_BLT_SEL A_PRE_N A_SEL_P<25> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<24> A_BLC<24> A_BLC_SEL A_BLT<24> A_BLT_SEL A_PRE_N A_SEL_P<24> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<23> A_BLC<23> A_BLC_SEL A_BLT<23> A_BLT_SEL A_PRE_N A_SEL_P<23> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<22> A_BLC<22> A_BLC_SEL A_BLT<22> A_BLT_SEL A_PRE_N A_SEL_P<22> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<21> A_BLC<21> A_BLC_SEL A_BLT<21> A_BLT_SEL A_PRE_N A_SEL_P<21> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<20> A_BLC<20> A_BLC_SEL A_BLT<20> A_BLT_SEL A_PRE_N A_SEL_P<20> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<19> A_BLC<19> A_BLC_SEL A_BLT<19> A_BLT_SEL A_PRE_N A_SEL_P<19> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<18> A_BLC<18> A_BLC_SEL A_BLT<18> A_BLT_SEL A_PRE_N A_SEL_P<18> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<17> A_BLC<17> A_BLC_SEL A_BLT<17> A_BLT_SEL A_PRE_N A_SEL_P<17> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<16> A_BLC<16> A_BLC_SEL A_BLT<16> A_BLT_SEL A_PRE_N A_SEL_P<16> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<15> A_BLC<15> A_BLC_SEL A_BLT<15> A_BLT_SEL A_PRE_N A_SEL_P<15> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<14> A_BLC<14> A_BLC_SEL A_BLT<14> A_BLT_SEL A_PRE_N A_SEL_P<14> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<13> A_BLC<13> A_BLC_SEL A_BLT<13> A_BLT_SEL A_PRE_N A_SEL_P<13> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<12> A_BLC<12> A_BLC_SEL A_BLT<12> A_BLT_SEL A_PRE_N A_SEL_P<12> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<11> A_BLC<11> A_BLC_SEL A_BLT<11> A_BLT_SEL A_PRE_N A_SEL_P<11> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<10> A_BLC<10> A_BLC_SEL A_BLT<10> A_BLT_SEL A_PRE_N A_SEL_P<10> 
+ A_WR_ONE A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<9> A_BLC<9> A_BLC_SEL A_BLT<9> A_BLT_SEL A_PRE_N A_SEL_P<9> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<8> A_BLC<8> A_BLC_SEL A_BLT<8> A_BLT_SEL A_PRE_N A_SEL_P<8> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<7> A_BLC<7> A_BLC_SEL A_BLT<7> A_BLT_SEL A_PRE_N A_SEL_P<7> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<6> A_BLC<6> A_BLC_SEL A_BLT<6> A_BLT_SEL A_PRE_N A_SEL_P<6> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<5> A_BLC<5> A_BLC_SEL A_BLT<5> A_BLT_SEL A_PRE_N A_SEL_P<5> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<4> A_BLC<4> A_BLC_SEL A_BLT<4> A_BLT_SEL A_PRE_N A_SEL_P<4> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<3> A_BLC<3> A_BLC_SEL A_BLT<3> A_BLT_SEL A_PRE_N A_SEL_P<3> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<2> A_BLC<2> A_BLC_SEL A_BLT<2> A_BLT_SEL A_PRE_N A_SEL_P<2> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<1> A_BLC<1> A_BLC_SEL A_BLT<1> A_BLT_SEL A_PRE_N A_SEL_P<1> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_BLTMUX<0> A_BLC<0> A_BLC_SEL A_BLT<0> A_BLT_SEL A_PRE_N A_SEL_P<0> A_WR_ONE 
+ A_WR_ZERO VDD VSS / RM_IHPSG13_2048x64_c2_1P_BLDRV
XA_CAPS<17> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<16> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<15> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<14> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<13> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<12> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<11> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<10> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<9> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<8> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<7> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<6> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX8
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X6
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X6
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<31> net23<0> A_SEL_P<31> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<30> net23<1> A_SEL_P<30> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<29> net23<2> A_SEL_P<29> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<28> net23<3> A_SEL_P<28> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<27> net23<4> A_SEL_P<27> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<26> net23<5> A_SEL_P<26> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<25> net23<6> A_SEL_P<25> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<24> net23<7> A_SEL_P<24> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<23> net23<8> A_SEL_P<23> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<22> net23<9> A_SEL_P<22> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<21> net23<10> A_SEL_P<21> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<20> net23<11> A_SEL_P<20> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<19> net23<12> A_SEL_P<19> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<18> net23<13> A_SEL_P<18> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<17> net23<14> A_SEL_P<17> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<16> net23<15> A_SEL_P<16> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<15> net23<16> A_SEL_P<15> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<14> net23<17> A_SEL_P<14> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<13> net23<18> A_SEL_P<13> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<12> net23<19> A_SEL_P<12> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<11> net23<20> A_SEL_P<11> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<10> net23<21> A_SEL_P<10> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<9> net23<22> A_SEL_P<9> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<8> net23<23> A_SEL_P<8> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<7> net23<24> A_SEL_P<7> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<6> net23<25> A_SEL_P<6> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<5> net23<26> A_SEL_P<5> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<4> net23<27> A_SEL_P<4> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<3> net23<28> A_SEL_P<3> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<2> net23<29> A_SEL_P<2> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<1> net23<30> A_SEL_P<1> VDD VSS / RSC_IHPSG13_INVX2
XA_DEC3INV<0> net23<31> A_SEL_P<0> VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net21 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_DEC3<31> A_P1<1> A_P0<1> A_ADDR_DEC<7> net23<0> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<30> A_P1<1> A_P0<1> A_ADDR_DEC<6> net23<1> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<29> A_P1<1> A_P0<1> A_ADDR_DEC<5> net23<2> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<28> A_P1<1> A_P0<1> A_ADDR_DEC<4> net23<3> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<27> A_P1<1> A_P0<1> A_ADDR_DEC<3> net23<4> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<26> A_P1<1> A_P0<1> A_ADDR_DEC<2> net23<5> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<25> A_P1<1> A_P0<1> A_ADDR_DEC<1> net23<6> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<24> A_P1<1> A_P0<1> A_ADDR_DEC<0> net23<7> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<23> A_P1<1> A_N0<1> A_ADDR_DEC<7> net23<8> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<22> A_P1<1> A_N0<1> A_ADDR_DEC<6> net23<9> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<21> A_P1<1> A_N0<1> A_ADDR_DEC<5> net23<10> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<20> A_P1<1> A_N0<1> A_ADDR_DEC<4> net23<11> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<19> A_P1<1> A_N0<1> A_ADDR_DEC<3> net23<12> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<18> A_P1<1> A_N0<1> A_ADDR_DEC<2> net23<13> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<17> A_P1<1> A_N0<1> A_ADDR_DEC<1> net23<14> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<16> A_P1<1> A_N0<1> A_ADDR_DEC<0> net23<15> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<15> A_N1<0> A_P0<0> A_ADDR_DEC<7> net23<16> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<14> A_N1<0> A_P0<0> A_ADDR_DEC<6> net23<17> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<13> A_N1<0> A_P0<0> A_ADDR_DEC<5> net23<18> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<12> A_N1<0> A_P0<0> A_ADDR_DEC<4> net23<19> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<11> A_N1<0> A_P0<0> A_ADDR_DEC<3> net23<20> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<10> A_N1<0> A_P0<0> A_ADDR_DEC<2> net23<21> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<9> A_N1<0> A_P0<0> A_ADDR_DEC<1> net23<22> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<8> A_N1<0> A_P0<0> A_ADDR_DEC<0> net23<23> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<7> A_N1<0> A_N0<0> A_ADDR_DEC<7> net23<24> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<6> A_N1<0> A_N0<0> A_ADDR_DEC<6> net23<25> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<5> A_N1<0> A_N0<0> A_ADDR_DEC<5> net23<26> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<4> A_N1<0> A_N0<0> A_ADDR_DEC<4> net23<27> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<3> A_N1<0> A_N0<0> A_ADDR_DEC<3> net23<28> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<2> A_N1<0> A_N0<0> A_ADDR_DEC<2> net23<29> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<1> A_N1<0> A_N0<0> A_ADDR_DEC<1> net23<30> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_DEC3<0> A_N1<0> A_N0<0> A_ADDR_DEC<0> net23<31> VDD VSS / 
+ RSC_IHPSG13_NAND3X2
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDRV13X12 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI1<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX12
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX12
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_WLDRV16X12 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX12
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX12
.ENDS



.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDRV13X8 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XI1<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RSC_IHPSG13_WLDRVX8 A Z VDD VSS
MN1 Z net6 VSS VSS nmos m=1 w=1.41u l=130.00n ng=2 nrd=0 nrs=0
MN0 net6 A VSS VSS nmos m=1 w=1.8u l=130.00n ng=2 nrd=0 nrs=0
MP1 Z net6 VDD VDD pmos m=1 w=6.48u l=130.00n ng=4 nrd=0 nrs=0
MP0 net6 A VDD VDD pmos m=1 w=900.0n l=130.00n ng=1 nrd=0 nrs=0
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_WLDRV16X8 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX8
.ENDS



.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDEC2 ACLK_N ADDR<1> ADDR<0> ADDR_COL<1> ADDR_COL<0> 
+ ADDR_DEC<7> ADDR_DEC<6> ADDR_DEC<5> ADDR_DEC<4> ADDR_DEC<3> ADDR_DEC<2> 
+ ADDR_DEC<1> ADDR_DEC<0> BIST_ADDR<1> BIST_ADDR<0> BIST_EN_I VDD VSS
XI16<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI16<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI18<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI1<3> PADR<0> PADR<1> addr_n<3> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<2> NADR<0> PADR<1> addr_n<2> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<1> PADR<0> NADR<1> addr_n<1> VDD VSS / RSC_IHPSG13_NAND2X2
XI1<0> NADR<0> NADR<1> addr_n<0> VDD VSS / RSC_IHPSG13_NAND2X2
XI17<1> ADDR_COL<1> VDD VSS / RSC_IHPSG13_TIEL
XI17<0> ADDR_COL<0> VDD VSS / RSC_IHPSG13_TIEL
XI14<3> ADDR_DEC<7> VDD VSS / RSC_IHPSG13_TIEL
XI14<2> ADDR_DEC<6> VDD VSS / RSC_IHPSG13_TIEL
XI14<1> ADDR_DEC<5> VDD VSS / RSC_IHPSG13_TIEL
XI14<0> ADDR_DEC<4> VDD VSS / RSC_IHPSG13_TIEL
XI13<1> NADR<1> PADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI13<0> NADR<0> PADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI3<1> padr_int<1> NADR<1> VDD VSS / RSC_IHPSG13_INVX2
XI3<0> padr_int<0> NADR<0> VDD VSS / RSC_IHPSG13_INVX2
XI2<3> addr_n<3> ADDR_DEC<3> VDD VSS / RSC_IHPSG13_INVX2
XI2<2> addr_n<2> ADDR_DEC<2> VDD VSS / RSC_IHPSG13_INVX2
XI2<1> addr_n<1> ADDR_DEC<1> VDD VSS / RSC_IHPSG13_INVX2
XI2<0> addr_n<0> ADDR_DEC<0> VDD VSS / RSC_IHPSG13_INVX2
XDFF<1> BIST_EN_I BIST_ADDR<1> ACLK_N ADDR<1> padr_int<1> net12<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR<0> ACLK_N ADDR<0> padr_int<0> net12<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI15<5> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI15<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI19<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLCTRL2 A_ADDR_DEC<3> A_ADDR_DEC<2> A_ADDR_DEC<1> 
+ A_ADDR_DEC<0> A_BIST_BM_I A_BIST_DW_I A_BIST_EN_I A_BLC<3> A_BLC<2> A_BLC<1> 
+ A_BLC<0> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_BM_I A_DCLK_B_L A_DCLK_B_R 
+ A_DCLK_L A_DCLK_R A_DR_O A_DW_I A_RCLK_B_L A_RCLK_B_R A_RCLK_L A_RCLK_R 
+ A_TIEH_O A_WCLK_B_L A_WCLK_B_R A_WCLK_L A_WCLK_R B_ADDR_DEC<3> B_ADDR_DEC<2> 
+ B_ADDR_DEC<1> B_ADDR_DEC<0> B_BIST_BM_I B_BIST_DW_I B_BIST_EN_I B_BLC<3> 
+ B_BLC<2> B_BLC<1> B_BLC<0> B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BM_I 
+ B_DCLK_B_L B_DCLK_B_R B_DCLK_L B_DCLK_R B_DR_O B_DW_I B_RCLK_B_L B_RCLK_B_R 
+ B_RCLK_L B_RCLK_R B_TIEH_O B_WCLK_B_L B_WCLK_B_R B_WCLK_L B_WCLK_R VDD 
+ VSS
XB_DREG B_BIST_EN_I B_BIST_DW_I B_DCLK_B_L B_DW_I B_DI_R net046 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XB_BREG B_BIST_EN_I B_BIST_BM_I B_DCLK_B_L B_BM_I B_BM_R net045 VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XA_DREG A_BIST_EN_I A_BIST_DW_I A_DCLK_B_L A_DW_I A_DI_R net22 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XA_BREG A_BIST_EN_I A_BIST_BM_I A_DCLK_B_L A_BM_I A_BM_R net23 VDD VSS 
+ / RSC_IHPSG13_DFNQMX2IX1
XB_CAPS VDD VSS / RSC_IHPSG13_FILLCAP4
XA_CAPS VDD VSS / RSC_IHPSG13_FILLCAP4
XB_I75 B_DI_R B_DO_WRITE_P B_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XB_I80 B_RCLK_B_L B_WCLK_B_L net041 VDD VSS / RSC_IHPSG13_AND2X2
XB_I76 B_DI_N B_DO_WRITE_P B_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XA_I80 A_RCLK_B_L A_WCLK_B_L net21 VDD VSS / RSC_IHPSG13_AND2X2
XA_I75 A_DI_R A_DO_WRITE_P A_WR_ONE VDD VSS / RSC_IHPSG13_AND2X2
XA_I76 A_DI_N A_DO_WRITE_P A_WR_ZERO VDD VSS / RSC_IHPSG13_AND2X2
XB_I44 B_WCLK_B_L B_BM_N B_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XA_I44 A_WCLK_B_L A_BM_N A_DO_WRITE_P VDD VSS / RSC_IHPSG13_NOR2X2
XB_I81 net041 B_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XA_I81 net21 A_PRE_N VDD VSS / RSC_IHPSG13_CINVX4_WN
XB_BM_TIEH B_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_BM_TIEH A_TIEH_O VDD VSS / RSC_IHPSG13_TIEH
XA_I89 A_DCLK_B_L A_DCLK_B_R / RSC_IHPSG13_MET3RES
XA_I88 A_DCLK_L A_DCLK_R / RSC_IHPSG13_MET3RES
XA_I87 A_WCLK_L A_WCLK_R / RSC_IHPSG13_MET3RES
XA_I91 A_RCLK_B_L A_RCLK_B_R / RSC_IHPSG13_MET3RES
XB_I87 B_WCLK_L B_WCLK_R / RSC_IHPSG13_MET3RES
XB_I88 B_DCLK_L B_DCLK_R / RSC_IHPSG13_MET3RES
XB_I89 B_DCLK_B_L B_DCLK_B_R / RSC_IHPSG13_MET3RES
XB_I90 B_WCLK_B_L B_WCLK_B_R / RSC_IHPSG13_MET3RES
XB_R2 B_RCLK_L B_RCLK_R / RSC_IHPSG13_MET3RES
XB_I91 B_RCLK_B_L B_RCLK_B_R / RSC_IHPSG13_MET3RES
XA_R2 A_RCLK_L A_RCLK_R / RSC_IHPSG13_MET3RES
XA_I90 A_WCLK_B_L A_WCLK_B_R / RSC_IHPSG13_MET3RES
XAB_BLMUX A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLC_SEL A_BLT<3> A_BLT<2> 
+ A_BLT<1> A_BLT<0> A_BLT_SEL A_PRE_N A_ADDR_DEC<3> A_ADDR_DEC<2> 
+ A_ADDR_DEC<1> A_ADDR_DEC<0> A_WR_ONE A_WR_ZERO B_BLC<3> B_BLC<2> B_BLC<1> 
+ B_BLC<0> B_BLC_SEL B_BLT<3> B_BLT<2> B_BLT<1> B_BLT<0> B_BLT_SEL B_PRE_N 
+ B_ADDR_DEC<3> B_ADDR_DEC<2> B_ADDR_DEC<1> B_ADDR_DEC<0> B_WR_ONE B_WR_ZERO 
+ VDD VSS / RM_IHPSG13_2048x64_c2_2P_BLDRV
XB_ISENSE B_SAE B_BLC_SEL B_BLT_SEL net039 net040 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XA_ISENSE A_SAE A_BLC_SEL A_BLT_SEL net19 net20 VDD VSS / 
+ RSC_IHPSG13_DFPQD_MSAFFX2
XB_I78 B_RCLK_B_L B_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XA_I78 A_RCLK_B_L A_SAE VDD VSS / RSC_IHPSG13_CBUFX2
XB_I83 B_BM_R B_BM_N VDD VSS / RSC_IHPSG13_INVX2
XB_I49 B_DI_R B_DI_N VDD VSS / RSC_IHPSG13_INVX2
XA_I83 A_BM_R A_BM_N VDD VSS / RSC_IHPSG13_INVX2
XA_I49 A_DI_R A_DI_N VDD VSS / RSC_IHPSG13_INVX2
XB_I51 net039 B_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I51 net19 A_DR_O VDD VSS / RSC_IHPSG13_INVX4
XA_I69 A_DCLK_L A_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_I50 A_WCLK_L A_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XA_EBUF A_RCLK_L A_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_EBUF B_RCLK_L B_RCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I50 B_WCLK_L B_WCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
XB_I69 B_DCLK_L B_DCLK_B_L VDD VSS / RSC_IHPSG13_CINVX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_COLDRV13_FILL4C2 VDD VSS
XI0<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWDEC7 ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> 
+ ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<127> WL_O<126> 
+ WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> 
+ WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> 
+ WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> WL_O<105> 
+ WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> WL_O<98> WL_O<97> 
+ WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> WL_O<90> WL_O<89> 
+ WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> WL_O<82> WL_O<81> 
+ WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> WL_O<74> WL_O<73> 
+ WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> WL_O<66> WL_O<65> 
+ WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> WL_O<58> WL_O<57> 
+ WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> WL_O<50> WL_O<49> 
+ WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> WL_O<42> WL_O<41> 
+ WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> WL_O<34> WL_O<33> 
+ WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> WL_O<26> WL_O<25> 
+ WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> WL_O<18> WL_O<17> 
+ WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC03
XDEC01<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC01
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC02
XDEC00<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_2P_DEC00
XI0 ADDR_N_I<7> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWREG7 ACLK_N_I ADDR_I<6> ADDR_I<5> ADDR_I<4> ADDR_I<3> 
+ ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<6> 
+ BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> 
+ BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<0> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWDEC4 ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> 
+ CS_I ECLK_I WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XSEL ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I ECLK_H<1> 
+ ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> 
+ WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> 
+ WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_2P_DEC04
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_2P_ROWREG4 ACLK_N_I ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net7<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net7<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net7<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net7<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI12<4> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<3> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<2> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI12<0> VDD VSS / RSC_IHPSG13_FILLCAP4
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_TAP BLC BLT NW PW VDD VSS
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_TAP A_BLC<1> A_BLC<0> A_BLT<1> A_BLT<0> 
+ VDD_CORE VSS
XITAP<1> A_BLC<1> A_BLT<1> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_1P_BITKIT_TAP
XITAP<0> A_BLC<0> A_BLT<0> VDD_CORE VSS VDD_CORE VSS 
+ / RM_IHPSG13_2048x64_c2_1P_BITKIT_TAP
XIEDGEBP_COL1<1> BLC<1> BLT<1> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL1<0> BLC<1> BLT<1> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL2<1> BLC<0> BLT<0> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB
XIEDGEBP_COL2<0> BLC<0> BLT<0> VDD_CORE VSS VDD_CORE 
+ VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_EDGE_TB
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_TAP_LR VDD_CORE VSS
XCORNER<1> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER
XCORNER<0> VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_CORNER
XTAP_BORDER VDD_CORE VSS VDD_CORE VSS / 
+ RM_IHPSG13_2048x64_c2_1P_BITKIT_TAP_LR
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_DEC03 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XI0 VDD VSS / RSC_IHPSG13_FILLCAP4
XDEC ADDR<1> ADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_DEC02 ADDR<1> ADDR<0> CS CS_OUT VDD VSS
XDECINV net1 CS_OUT VDD VSS / RSC_IHPSG13_INVX4
XDEC ADDR<1> NADDR<0> CS net1 VDD VSS / RSC_IHPSG13_NAND3X2
XI2 VDD VSS / RSC_IHPSG13_FILLCAP4
XADDRINV ADDR<0> NADDR<0> VDD VSS / RSC_IHPSG13_INVX2
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWDEC8 ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> 
+ ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<255> 
+ WL_O<254> WL_O<253> WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> 
+ WL_O<247> WL_O<246> WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> 
+ WL_O<240> WL_O<239> WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> 
+ WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> 
+ WL_O<226> WL_O<225> WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> 
+ WL_O<205> WL_O<204> WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> 
+ WL_O<198> WL_O<197> WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> 
+ WL_O<191> WL_O<190> WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> 
+ WL_O<184> WL_O<183> WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> 
+ WL_O<177> WL_O<176> WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> 
+ WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> 
+ WL_O<163> WL_O<162> WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> 
+ WL_O<156> WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> 
+ WL_O<149> WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> 
+ WL_O<142> WL_O<141> WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> 
+ WL_O<135> WL_O<134> WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> 
+ WL_O<128> WL_O<127> WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> 
+ WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> 
+ WL_O<114> WL_O<113> WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> 
+ WL_O<92> WL_O<91> WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> 
+ WL_O<84> WL_O<83> WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> 
+ WL_O<76> WL_O<75> WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> 
+ WL_O<68> WL_O<67> WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> 
+ WL_O<60> WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> 
+ WL_O<52> WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> 
+ WL_O<44> WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> 
+ WL_O<36> WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> 
+ WL_O<28> WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> 
+ WL_O<20> WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> 
+ WL_O<12> WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> 
+ WL_O<3> WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC10<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC00<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XDEC01<4> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS04<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS04<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWREG8 ACLK_N_I ADDR_I<7> ADDR_I<6> ADDR_I<5> ADDR_I<4> 
+ ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<7> ADDR_N_O<6> ADDR_N_O<5> 
+ ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<7> 
+ BIST_ADDR_I<6> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> 
+ BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWDEC9 ADDR_N_I<8> ADDR_N_I<7> ADDR_N_I<6> ADDR_N_I<5> 
+ ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I 
+ WL_O<511> WL_O<510> WL_O<509> WL_O<508> WL_O<507> WL_O<506> WL_O<505> 
+ WL_O<504> WL_O<503> WL_O<502> WL_O<501> WL_O<500> WL_O<499> WL_O<498> 
+ WL_O<497> WL_O<496> WL_O<495> WL_O<494> WL_O<493> WL_O<492> WL_O<491> 
+ WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> WL_O<484> 
+ WL_O<483> WL_O<482> WL_O<481> WL_O<480> WL_O<479> WL_O<478> WL_O<477> 
+ WL_O<476> WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> 
+ WL_O<469> WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> WL_O<463> 
+ WL_O<462> WL_O<461> WL_O<460> WL_O<459> WL_O<458> WL_O<457> WL_O<456> 
+ WL_O<455> WL_O<454> WL_O<453> WL_O<452> WL_O<451> WL_O<450> WL_O<449> 
+ WL_O<448> WL_O<447> WL_O<446> WL_O<445> WL_O<444> WL_O<443> WL_O<442> 
+ WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> WL_O<436> WL_O<435> 
+ WL_O<434> WL_O<433> WL_O<432> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> WL_O<415> WL_O<414> 
+ WL_O<413> WL_O<412> WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> 
+ WL_O<406> WL_O<405> WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> 
+ WL_O<399> WL_O<398> WL_O<397> WL_O<396> WL_O<395> WL_O<394> WL_O<393> 
+ WL_O<392> WL_O<391> WL_O<390> WL_O<389> WL_O<388> WL_O<387> WL_O<386> 
+ WL_O<385> WL_O<384> WL_O<383> WL_O<382> WL_O<381> WL_O<380> WL_O<379> 
+ WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> WL_O<372> 
+ WL_O<371> WL_O<370> WL_O<369> WL_O<368> WL_O<367> WL_O<366> WL_O<365> 
+ WL_O<364> WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> 
+ WL_O<357> WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> WL_O<351> 
+ WL_O<350> WL_O<349> WL_O<348> WL_O<347> WL_O<346> WL_O<345> WL_O<344> 
+ WL_O<343> WL_O<342> WL_O<341> WL_O<340> WL_O<339> WL_O<338> WL_O<337> 
+ WL_O<336> WL_O<335> WL_O<334> WL_O<333> WL_O<332> WL_O<331> WL_O<330> 
+ WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> WL_O<324> WL_O<323> 
+ WL_O<322> WL_O<321> WL_O<320> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> WL_O<303> WL_O<302> 
+ WL_O<301> WL_O<300> WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> 
+ WL_O<294> WL_O<293> WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> 
+ WL_O<287> WL_O<286> WL_O<285> WL_O<284> WL_O<283> WL_O<282> WL_O<281> 
+ WL_O<280> WL_O<279> WL_O<278> WL_O<277> WL_O<276> WL_O<275> WL_O<274> 
+ WL_O<273> WL_O<272> WL_O<271> WL_O<270> WL_O<269> WL_O<268> WL_O<267> 
+ WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> WL_O<260> 
+ WL_O<259> WL_O<258> WL_O<257> WL_O<256> WL_O<255> WL_O<254> WL_O<253> 
+ WL_O<252> WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> 
+ WL_O<245> WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> WL_O<239> 
+ WL_O<238> WL_O<237> WL_O<236> WL_O<235> WL_O<234> WL_O<233> WL_O<232> 
+ WL_O<231> WL_O<230> WL_O<229> WL_O<228> WL_O<227> WL_O<226> WL_O<225> 
+ WL_O<224> WL_O<223> WL_O<222> WL_O<221> WL_O<220> WL_O<219> WL_O<218> 
+ WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> WL_O<212> WL_O<211> 
+ WL_O<210> WL_O<209> WL_O<208> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> WL_O<191> WL_O<190> 
+ WL_O<189> WL_O<188> WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> 
+ WL_O<182> WL_O<181> WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> 
+ WL_O<175> WL_O<174> WL_O<173> WL_O<172> WL_O<171> WL_O<170> WL_O<169> 
+ WL_O<168> WL_O<167> WL_O<166> WL_O<165> WL_O<164> WL_O<163> WL_O<162> 
+ WL_O<161> WL_O<160> WL_O<159> WL_O<158> WL_O<157> WL_O<156> WL_O<155> 
+ WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> WL_O<148> 
+ WL_O<147> WL_O<146> WL_O<145> WL_O<144> WL_O<143> WL_O<142> WL_O<141> 
+ WL_O<140> WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> 
+ WL_O<133> WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> WL_O<127> 
+ WL_O<126> WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> 
+ WL_O<119> WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> 
+ WL_O<112> WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> 
+ WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> 
+ WL_O<98> WL_O<97> WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS
XL2<172> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<171> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<170> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<169> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<168> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<167> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<166> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<165> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<164> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<163> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<162> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<161> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<160> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<159> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<158> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<157> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<156> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<155> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<154> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<153> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<152> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<151> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<150> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<149> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<148> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<147> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<146> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<145> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<144> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<143> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<142> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<141> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<140> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<139> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<138> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<137> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<136> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<135> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<134> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<133> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<132> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<131> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<130> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<129> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<128> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<127> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<126> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<125> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<124> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<123> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<122> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<121> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<120> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<119> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<118> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<117> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<116> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<115> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<114> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<113> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<112> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<111> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<110> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<109> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<108> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<107> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<106> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<105> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<104> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<103> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<102> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<101> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<100> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<99> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<98> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<97> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<96> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<95> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<94> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<93> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<92> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<91> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<90> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<89> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<88> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<87> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<86> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<85> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<84> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<83> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<82> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<81> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<80> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<79> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<78> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<77> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<76> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<75> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<74> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<73> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<72> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<71> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<70> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<69> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<68> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<67> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<66> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<65> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<64> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<63> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<62> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<61> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<60> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<59> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<58> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<57> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<56> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<55> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<54> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<53> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<52> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<51> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<50> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<49> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<48> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<47> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<46> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<45> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XDEC11<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<31> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<27> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<23> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<19> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<15> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<11> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC00<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<28> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<24> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<20> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<16> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<12> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<8> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XSEL<31> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<31> ECLK_H<31> 
+ ECLK_H<32> ECLK_B<31> ECLK_B<32> WL_O<511> WL_O<510> WL_O<509> WL_O<508> 
+ WL_O<507> WL_O<506> WL_O<505> WL_O<504> WL_O<503> WL_O<502> WL_O<501> 
+ WL_O<500> WL_O<499> WL_O<498> WL_O<497> WL_O<496> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<30> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<30> ECLK_H<30> 
+ ECLK_H<31> ECLK_B<30> ECLK_B<31> WL_O<495> WL_O<494> WL_O<493> WL_O<492> 
+ WL_O<491> WL_O<490> WL_O<489> WL_O<488> WL_O<487> WL_O<486> WL_O<485> 
+ WL_O<484> WL_O<483> WL_O<482> WL_O<481> WL_O<480> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<29> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<29> ECLK_H<29> 
+ ECLK_H<30> ECLK_B<29> ECLK_B<30> WL_O<479> WL_O<478> WL_O<477> WL_O<476> 
+ WL_O<475> WL_O<474> WL_O<473> WL_O<472> WL_O<471> WL_O<470> WL_O<469> 
+ WL_O<468> WL_O<467> WL_O<466> WL_O<465> WL_O<464> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<28> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<28> ECLK_H<28> 
+ ECLK_H<29> ECLK_B<28> ECLK_B<29> WL_O<463> WL_O<462> WL_O<461> WL_O<460> 
+ WL_O<459> WL_O<458> WL_O<457> WL_O<456> WL_O<455> WL_O<454> WL_O<453> 
+ WL_O<452> WL_O<451> WL_O<450> WL_O<449> WL_O<448> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<27> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<27> ECLK_H<27> 
+ ECLK_H<28> ECLK_B<27> ECLK_B<28> WL_O<447> WL_O<446> WL_O<445> WL_O<444> 
+ WL_O<443> WL_O<442> WL_O<441> WL_O<440> WL_O<439> WL_O<438> WL_O<437> 
+ WL_O<436> WL_O<435> WL_O<434> WL_O<433> WL_O<432> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<26> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<26> ECLK_H<26> 
+ ECLK_H<27> ECLK_B<26> ECLK_B<27> WL_O<431> WL_O<430> WL_O<429> WL_O<428> 
+ WL_O<427> WL_O<426> WL_O<425> WL_O<424> WL_O<423> WL_O<422> WL_O<421> 
+ WL_O<420> WL_O<419> WL_O<418> WL_O<417> WL_O<416> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<25> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<25> ECLK_H<25> 
+ ECLK_H<26> ECLK_B<25> ECLK_B<26> WL_O<415> WL_O<414> WL_O<413> WL_O<412> 
+ WL_O<411> WL_O<410> WL_O<409> WL_O<408> WL_O<407> WL_O<406> WL_O<405> 
+ WL_O<404> WL_O<403> WL_O<402> WL_O<401> WL_O<400> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<24> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<24> ECLK_H<24> 
+ ECLK_H<25> ECLK_B<24> ECLK_B<25> WL_O<399> WL_O<398> WL_O<397> WL_O<396> 
+ WL_O<395> WL_O<394> WL_O<393> WL_O<392> WL_O<391> WL_O<390> WL_O<389> 
+ WL_O<388> WL_O<387> WL_O<386> WL_O<385> WL_O<384> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<23> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<23> ECLK_H<23> 
+ ECLK_H<24> ECLK_B<23> ECLK_B<24> WL_O<383> WL_O<382> WL_O<381> WL_O<380> 
+ WL_O<379> WL_O<378> WL_O<377> WL_O<376> WL_O<375> WL_O<374> WL_O<373> 
+ WL_O<372> WL_O<371> WL_O<370> WL_O<369> WL_O<368> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<22> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<22> ECLK_H<22> 
+ ECLK_H<23> ECLK_B<22> ECLK_B<23> WL_O<367> WL_O<366> WL_O<365> WL_O<364> 
+ WL_O<363> WL_O<362> WL_O<361> WL_O<360> WL_O<359> WL_O<358> WL_O<357> 
+ WL_O<356> WL_O<355> WL_O<354> WL_O<353> WL_O<352> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<21> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<21> ECLK_H<21> 
+ ECLK_H<22> ECLK_B<21> ECLK_B<22> WL_O<351> WL_O<350> WL_O<349> WL_O<348> 
+ WL_O<347> WL_O<346> WL_O<345> WL_O<344> WL_O<343> WL_O<342> WL_O<341> 
+ WL_O<340> WL_O<339> WL_O<338> WL_O<337> WL_O<336> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<20> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<20> ECLK_H<20> 
+ ECLK_H<21> ECLK_B<20> ECLK_B<21> WL_O<335> WL_O<334> WL_O<333> WL_O<332> 
+ WL_O<331> WL_O<330> WL_O<329> WL_O<328> WL_O<327> WL_O<326> WL_O<325> 
+ WL_O<324> WL_O<323> WL_O<322> WL_O<321> WL_O<320> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<19> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<19> ECLK_H<19> 
+ ECLK_H<20> ECLK_B<19> ECLK_B<20> WL_O<319> WL_O<318> WL_O<317> WL_O<316> 
+ WL_O<315> WL_O<314> WL_O<313> WL_O<312> WL_O<311> WL_O<310> WL_O<309> 
+ WL_O<308> WL_O<307> WL_O<306> WL_O<305> WL_O<304> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<18> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<18> ECLK_H<18> 
+ ECLK_H<19> ECLK_B<18> ECLK_B<19> WL_O<303> WL_O<302> WL_O<301> WL_O<300> 
+ WL_O<299> WL_O<298> WL_O<297> WL_O<296> WL_O<295> WL_O<294> WL_O<293> 
+ WL_O<292> WL_O<291> WL_O<290> WL_O<289> WL_O<288> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<17> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<17> ECLK_H<17> 
+ ECLK_H<18> ECLK_B<17> ECLK_B<18> WL_O<287> WL_O<286> WL_O<285> WL_O<284> 
+ WL_O<283> WL_O<282> WL_O<281> WL_O<280> WL_O<279> WL_O<278> WL_O<277> 
+ WL_O<276> WL_O<275> WL_O<274> WL_O<273> WL_O<272> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<16> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<16> ECLK_H<16> 
+ ECLK_H<17> ECLK_B<16> ECLK_B<17> WL_O<271> WL_O<270> WL_O<269> WL_O<268> 
+ WL_O<267> WL_O<266> WL_O<265> WL_O<264> WL_O<263> WL_O<262> WL_O<261> 
+ WL_O<260> WL_O<259> WL_O<258> WL_O<257> WL_O<256> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<15> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<15> ECLK_H<15> 
+ ECLK_H<16> ECLK_B<15> ECLK_B<16> WL_O<255> WL_O<254> WL_O<253> WL_O<252> 
+ WL_O<251> WL_O<250> WL_O<249> WL_O<248> WL_O<247> WL_O<246> WL_O<245> 
+ WL_O<244> WL_O<243> WL_O<242> WL_O<241> WL_O<240> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<14> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<14> ECLK_H<14> 
+ ECLK_H<15> ECLK_B<14> ECLK_B<15> WL_O<239> WL_O<238> WL_O<237> WL_O<236> 
+ WL_O<235> WL_O<234> WL_O<233> WL_O<232> WL_O<231> WL_O<230> WL_O<229> 
+ WL_O<228> WL_O<227> WL_O<226> WL_O<225> WL_O<224> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<13> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<13> ECLK_H<13> 
+ ECLK_H<14> ECLK_B<13> ECLK_B<14> WL_O<223> WL_O<222> WL_O<221> WL_O<220> 
+ WL_O<219> WL_O<218> WL_O<217> WL_O<216> WL_O<215> WL_O<214> WL_O<213> 
+ WL_O<212> WL_O<211> WL_O<210> WL_O<209> WL_O<208> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<12> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<12> ECLK_H<12> 
+ ECLK_H<13> ECLK_B<12> ECLK_B<13> WL_O<207> WL_O<206> WL_O<205> WL_O<204> 
+ WL_O<203> WL_O<202> WL_O<201> WL_O<200> WL_O<199> WL_O<198> WL_O<197> 
+ WL_O<196> WL_O<195> WL_O<194> WL_O<193> WL_O<192> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<11> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<11> ECLK_H<11> 
+ ECLK_H<12> ECLK_B<11> ECLK_B<12> WL_O<191> WL_O<190> WL_O<189> WL_O<188> 
+ WL_O<187> WL_O<186> WL_O<185> WL_O<184> WL_O<183> WL_O<182> WL_O<181> 
+ WL_O<180> WL_O<179> WL_O<178> WL_O<177> WL_O<176> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<10> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<10> ECLK_H<10> 
+ ECLK_H<11> ECLK_B<10> ECLK_B<11> WL_O<175> WL_O<174> WL_O<173> WL_O<172> 
+ WL_O<171> WL_O<170> WL_O<169> WL_O<168> WL_O<167> WL_O<166> WL_O<165> 
+ WL_O<164> WL_O<163> WL_O<162> WL_O<161> WL_O<160> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<9> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<9> ECLK_H<9> 
+ ECLK_H<10> ECLK_B<9> ECLK_B<10> WL_O<159> WL_O<158> WL_O<157> WL_O<156> 
+ WL_O<155> WL_O<154> WL_O<153> WL_O<152> WL_O<151> WL_O<150> WL_O<149> 
+ WL_O<148> WL_O<147> WL_O<146> WL_O<145> WL_O<144> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<8> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<8> ECLK_H<8> 
+ ECLK_H<9> ECLK_B<8> ECLK_B<9> WL_O<143> WL_O<142> WL_O<141> WL_O<140> 
+ WL_O<139> WL_O<138> WL_O<137> WL_O<136> WL_O<135> WL_O<134> WL_O<133> 
+ WL_O<132> WL_O<131> WL_O<130> WL_O<129> WL_O<128> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XDEC01<10> ADDR_N_I<9> ADDR_N_I<8> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<29> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<25> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<21> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<17> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<13> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<9> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC10<9> ADDR_N_I<7> ADDR_N_I<6> CS04<1> CS02<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<8> ADDR_N_I<7> ADDR_N_I<6> CS04<0> CS02<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<7> ADDR_N_I<5> ADDR_N_I<4> CS02<7> CS00<30> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<6> ADDR_N_I<5> ADDR_N_I<4> CS02<6> CS00<26> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<5> ADDR_N_I<5> ADDR_N_I<4> CS02<5> CS00<22> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<4> ADDR_N_I<5> ADDR_N_I<4> CS02<4> CS00<18> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<3> ADDR_N_I<5> ADDR_N_I<4> CS02<3> CS00<14> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<2> ADDR_N_I<5> ADDR_N_I<4> CS02<2> CS00<10> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS02<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS02<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XI0 ADDR_N_I<9> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWREG9 ACLK_N_I ADDR_I<8> ADDR_I<7> ADDR_I<6> ADDR_I<5> 
+ ADDR_I<4> ADDR_I<3> ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<8> ADDR_N_O<7> 
+ ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> 
+ ADDR_N_O<0> BIST_ADDR_I<8> BIST_ADDR_I<7> BIST_ADDR_I<6> BIST_ADDR_I<5> 
+ BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> 
+ BIST_EN_I VDD VSS
XINV<8> q_int<8> qn_int<8> VDD VSS / RSC_IHPSG13_CINVX2
XINV<7> q_int<7> qn_int<7> VDD VSS / RSC_IHPSG13_CINVX2
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<8> qn_int<8> ADDR_N_O<8> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<7> qn_int<7> ADDR_N_O<7> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<8> BIST_EN_I BIST_ADDR_I<8> ACLK_N_I ADDR_I<8> q_int<8> net04<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<7> BIST_EN_I BIST_ADDR_I<7> ACLK_N_I ADDR_I<7> q_int<7> net04<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net04<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net04<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net04<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net04<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net04<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net04<7> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net04<8> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWDEC7 ADDR_N_I<6> ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> 
+ ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<127> WL_O<126> 
+ WL_O<125> WL_O<124> WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> 
+ WL_O<118> WL_O<117> WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> 
+ WL_O<111> WL_O<110> WL_O<109> WL_O<108> WL_O<107> WL_O<106> WL_O<105> 
+ WL_O<104> WL_O<103> WL_O<102> WL_O<101> WL_O<100> WL_O<99> WL_O<98> WL_O<97> 
+ WL_O<96> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> WL_O<90> WL_O<89> 
+ WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> WL_O<82> WL_O<81> 
+ WL_O<80> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> WL_O<74> WL_O<73> 
+ WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> WL_O<66> WL_O<65> 
+ WL_O<64> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> WL_O<58> WL_O<57> 
+ WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> WL_O<50> WL_O<49> 
+ WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> WL_O<42> WL_O<41> 
+ WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> WL_O<34> WL_O<33> 
+ WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> WL_O<26> WL_O<25> 
+ WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> WL_O<18> WL_O<17> 
+ WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> WL_O<10> WL_O<9> 
+ WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> WL_O<1> WL_O<0> 
+ VDD VSS
XDEC11<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<7> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC11<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC10<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<6> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XDEC10<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XSEL<7> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<7> ECLK_H<7> 
+ ECLK_H<8> ECLK_B<7> ECLK_B<8> WL_O<127> WL_O<126> WL_O<125> WL_O<124> 
+ WL_O<123> WL_O<122> WL_O<121> WL_O<120> WL_O<119> WL_O<118> WL_O<117> 
+ WL_O<116> WL_O<115> WL_O<114> WL_O<113> WL_O<112> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<6> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<6> ECLK_H<6> 
+ ECLK_H<7> ECLK_B<6> ECLK_B<7> WL_O<111> WL_O<110> WL_O<109> WL_O<108> 
+ WL_O<107> WL_O<106> WL_O<105> WL_O<104> WL_O<103> WL_O<102> WL_O<101> 
+ WL_O<100> WL_O<99> WL_O<98> WL_O<97> WL_O<96> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<5> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<5> ECLK_H<5> 
+ ECLK_H<6> ECLK_B<5> ECLK_B<6> WL_O<95> WL_O<94> WL_O<93> WL_O<92> WL_O<91> 
+ WL_O<90> WL_O<89> WL_O<88> WL_O<87> WL_O<86> WL_O<85> WL_O<84> WL_O<83> 
+ WL_O<82> WL_O<81> WL_O<80> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<4> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<4> ECLK_H<4> 
+ ECLK_H<5> ECLK_B<4> ECLK_B<5> WL_O<79> WL_O<78> WL_O<77> WL_O<76> WL_O<75> 
+ WL_O<74> WL_O<73> WL_O<72> WL_O<71> WL_O<70> WL_O<69> WL_O<68> WL_O<67> 
+ WL_O<66> WL_O<65> WL_O<64> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XDEC00<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<4> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC00<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC01<2> ADDR_N_I<7> ADDR_N_I<6> CS_I CS04<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<1> ADDR_N_I<5> ADDR_N_I<4> CS04<1> CS00<5> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC01<0> ADDR_N_I<5> ADDR_N_I<4> CS04<0> CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XL2<44> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<43> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<42> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<41> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<40> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<39> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<38> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<37> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<36> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<35> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<34> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<33> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<32> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<31> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<30> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<29> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<28> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<27> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<26> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<25> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
XI0 ADDR_N_I<7> VDD VSS / RSC_IHPSG13_TIEL
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWREG7 ACLK_N_I ADDR_I<6> ADDR_I<5> ADDR_I<4> ADDR_I<3> 
+ ADDR_I<2> ADDR_I<1> ADDR_I<0> ADDR_N_O<6> ADDR_N_O<5> ADDR_N_O<4> 
+ ADDR_N_O<3> ADDR_N_O<2> ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<6> 
+ BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> BIST_ADDR_I<2> BIST_ADDR_I<1> 
+ BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<6> q_int<6> qn_int<6> VDD VSS / RSC_IHPSG13_CINVX2
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<6> qn_int<6> ADDR_N_O<6> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<6> BIST_EN_I BIST_ADDR_I<6> ACLK_N_I ADDR_I<6> q_int<6> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<6> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS

.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLDRV13X8 ADDR_COL_I<1> ADDR_COL_I<0> ADDR_COL_O<1> 
+ ADDR_COL_O<0> ADDR_DEC_I<7> ADDR_DEC_I<6> ADDR_DEC_I<5> ADDR_DEC_I<4> 
+ ADDR_DEC_I<3> ADDR_DEC_I<2> ADDR_DEC_I<1> ADDR_DEC_I<0> ADDR_DEC_O<7> 
+ ADDR_DEC_O<6> ADDR_DEC_O<5> ADDR_DEC_O<4> ADDR_DEC_O<3> ADDR_DEC_O<2> 
+ ADDR_DEC_O<1> ADDR_DEC_O<0> DCLK_I DCLK_O RCLK_I RCLK_O WCLK_I WCLK_O 
+ VDD VSS
XI0<1> VDD VSS / RSC_IHPSG13_FILLCAP4
XI0<0> VDD VSS / RSC_IHPSG13_FILLCAP4
XADDR_COL_DRV<1> ADDR_COL_I<1> ADDR_COL_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_COL_DRV<0> ADDR_COL_I<0> ADDR_COL_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<7> ADDR_DEC_I<7> ADDR_DEC_O<7> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<6> ADDR_DEC_I<6> ADDR_DEC_O<6> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<5> ADDR_DEC_I<5> ADDR_DEC_O<5> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<4> ADDR_DEC_I<4> ADDR_DEC_O<4> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<3> ADDR_DEC_I<3> ADDR_DEC_O<3> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<2> ADDR_DEC_I<2> ADDR_DEC_O<2> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<1> ADDR_DEC_I<1> ADDR_DEC_O<1> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XADDR_DEC_DRV<0> ADDR_DEC_I<0> ADDR_DEC_O<0> VDD VSS / 
+ RSC_IHPSG13_CBUFX8
XDCLK_DRV DCLK_I DCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XRCLK_DRV RCLK_I RCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
XWCLK_DRV WCLK_I WCLK_O VDD VSS / RSC_IHPSG13_CBUFX8
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_WLDRV16X8 A<15> A<14> A<13> A<12> A<11> A<10> A<9> A<8> 
+ A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> Z<15> Z<14> Z<13> Z<12> Z<11> Z<10> 
+ Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> VDD VSS
XBUF<15> A<15> Z<15> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<14> A<14> Z<14> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<13> A<13> Z<13> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<12> A<12> Z<12> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<11> A<11> Z<11> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<10> A<10> Z<10> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<9> A<9> Z<9> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<8> A<8> Z<8> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<7> A<7> Z<7> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<6> A<6> Z<6> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<5> A<5> Z<5> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<4> A<4> Z<4> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<3> A<3> Z<3> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<2> A<2> Z<2> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<1> A<1> Z<1> VDD VSS / RSC_IHPSG13_WLDRVX8
XBUF<0> A<0> Z<0> VDD VSS / RSC_IHPSG13_WLDRVX8
.ENDS



.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWDEC6 ADDR_N_I<5> ADDR_N_I<4> ADDR_N_I<3> ADDR_N_I<2> 
+ ADDR_N_I<1> ADDR_N_I<0> CS_I ECLK_I WL_O<63> WL_O<62> WL_O<61> WL_O<60> 
+ WL_O<59> WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> 
+ WL_O<51> WL_O<50> WL_O<49> WL_O<48> WL_O<47> WL_O<46> WL_O<45> WL_O<44> 
+ WL_O<43> WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> 
+ WL_O<35> WL_O<34> WL_O<33> WL_O<32> WL_O<31> WL_O<30> WL_O<29> WL_O<28> 
+ WL_O<27> WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> 
+ WL_O<19> WL_O<18> WL_O<17> WL_O<16> WL_O<15> WL_O<14> WL_O<13> WL_O<12> 
+ WL_O<11> WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> 
+ WL_O<2> WL_O<1> WL_O<0> VDD VSS
XDEC11 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<3> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC03
XDEC00 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<0> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC00
XDEC01 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<1> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC01
XDEC10 ADDR_N_I<5> ADDR_N_I<4> CS_I CS00<2> VDD VSS / 
+ RM_IHPSG13_2048x64_c2_1P_DEC02
XSEL<3> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<3> ECLK_H<3> 
+ ECLK_H<4> ECLK_B<3> ECLK_B<4> WL_O<63> WL_O<62> WL_O<61> WL_O<60> WL_O<59> 
+ WL_O<58> WL_O<57> WL_O<56> WL_O<55> WL_O<54> WL_O<53> WL_O<52> WL_O<51> 
+ WL_O<50> WL_O<49> WL_O<48> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<2> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<2> ECLK_H<2> 
+ ECLK_H<3> ECLK_B<2> ECLK_B<3> WL_O<47> WL_O<46> WL_O<45> WL_O<44> WL_O<43> 
+ WL_O<42> WL_O<41> WL_O<40> WL_O<39> WL_O<38> WL_O<37> WL_O<36> WL_O<35> 
+ WL_O<34> WL_O<33> WL_O<32> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<1> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<1> ECLK_H<1> 
+ ECLK_H<2> ECLK_B<1> ECLK_B<2> WL_O<31> WL_O<30> WL_O<29> WL_O<28> WL_O<27> 
+ WL_O<26> WL_O<25> WL_O<24> WL_O<23> WL_O<22> WL_O<21> WL_O<20> WL_O<19> 
+ WL_O<18> WL_O<17> WL_O<16> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XSEL<0> ADDR_N_I<3> ADDR_N_I<2> ADDR_N_I<1> ADDR_N_I<0> CS00<0> ECLK_I 
+ ECLK_H<1> ECLK_B<0> ECLK_B<1> WL_O<15> WL_O<14> WL_O<13> WL_O<12> WL_O<11> 
+ WL_O<10> WL_O<9> WL_O<8> WL_O<7> WL_O<6> WL_O<5> WL_O<4> WL_O<3> WL_O<2> 
+ WL_O<1> WL_O<0> VDD VSS / RM_IHPSG13_2048x64_c2_1P_DEC04
XL2<24> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<23> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<22> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<21> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<20> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<19> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<18> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<17> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<16> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<15> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<14> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<13> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XL2<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS
.SUBCKT RM_IHPSG13_2048x64_c2_1P_ROWREG6 ACLK_N_I ADDR_I<5> ADDR_I<4> ADDR_I<3> ADDR_I<2> 
+ ADDR_I<1> ADDR_I<0> ADDR_N_O<5> ADDR_N_O<4> ADDR_N_O<3> ADDR_N_O<2> 
+ ADDR_N_O<1> ADDR_N_O<0> BIST_ADDR_I<5> BIST_ADDR_I<4> BIST_ADDR_I<3> 
+ BIST_ADDR_I<2> BIST_ADDR_I<1> BIST_ADDR_I<0> BIST_EN_I VDD VSS
XINV<5> q_int<5> qn_int<5> VDD VSS / RSC_IHPSG13_CINVX2
XINV<4> q_int<4> qn_int<4> VDD VSS / RSC_IHPSG13_CINVX2
XINV<3> q_int<3> qn_int<3> VDD VSS / RSC_IHPSG13_CINVX2
XINV<2> q_int<2> qn_int<2> VDD VSS / RSC_IHPSG13_CINVX2
XINV<1> q_int<1> qn_int<1> VDD VSS / RSC_IHPSG13_CINVX2
XINV<0> q_int<0> qn_int<0> VDD VSS / RSC_IHPSG13_CINVX2
XDRV<5> qn_int<5> ADDR_N_O<5> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<4> qn_int<4> ADDR_N_O<4> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<3> qn_int<3> ADDR_N_O<3> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<2> qn_int<2> ADDR_N_O<2> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<1> qn_int<1> ADDR_N_O<1> VDD VSS / RSC_IHPSG13_CINVX8
XDRV<0> qn_int<0> ADDR_N_O<0> VDD VSS / RSC_IHPSG13_CINVX8
XDFF<5> BIST_EN_I BIST_ADDR_I<5> ACLK_N_I ADDR_I<5> q_int<5> net2<0> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<4> BIST_EN_I BIST_ADDR_I<4> ACLK_N_I ADDR_I<4> q_int<4> net2<1> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<3> BIST_EN_I BIST_ADDR_I<3> ACLK_N_I ADDR_I<3> q_int<3> net2<2> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<2> BIST_EN_I BIST_ADDR_I<2> ACLK_N_I ADDR_I<2> q_int<2> net2<3> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<1> BIST_EN_I BIST_ADDR_I<1> ACLK_N_I ADDR_I<1> q_int<1> net2<4> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XDFF<0> BIST_EN_I BIST_ADDR_I<0> ACLK_N_I ADDR_I<0> q_int<0> net2<5> VDD 
+ VSS / RSC_IHPSG13_DFNQMX2IX1
XI11<12> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<11> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<10> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<9> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<8> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<7> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<6> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<5> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<4> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<3> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<2> VDD VSS / RSC_IHPSG13_FILLCAP8
XI11<1> VDD VSS / RSC_IHPSG13_FILLCAP8
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0 A_BLC_BOT<1> A_BLC_BOT<0> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<511> A_LWL<510> A_LWL<509> A_LWL<508> A_LWL<507> A_LWL<506> A_LWL<505> A_LWL<504> A_LWL<503> A_LWL<502> A_LWL<501> A_LWL<500> A_LWL<499> A_LWL<498> A_LWL<497> A_LWL<496> A_LWL<495> A_LWL<494> A_LWL<493> A_LWL<492> A_LWL<491> A_LWL<490> A_LWL<489> A_LWL<488> A_LWL<487> A_LWL<486> A_LWL<485> A_LWL<484> A_LWL<483> A_LWL<482> A_LWL<481> A_LWL<480> A_LWL<479> A_LWL<478> A_LWL<477> A_LWL<476> A_LWL<475> A_LWL<474> A_LWL<473> A_LWL<472> A_LWL<471> A_LWL<470> A_LWL<469> A_LWL<468> A_LWL<467> A_LWL<466> A_LWL<465> A_LWL<464> A_LWL<463> A_LWL<462> A_LWL<461> A_LWL<460> A_LWL<459> A_LWL<458> A_LWL<457> A_LWL<456> A_LWL<455> A_LWL<454> A_LWL<453> A_LWL<452> A_LWL<451> A_LWL<450> A_LWL<449> A_LWL<448> A_LWL<447> A_LWL<446> A_LWL<445> A_LWL<444> A_LWL<443> A_LWL<442> A_LWL<441> A_LWL<440> A_LWL<439> A_LWL<438> A_LWL<437> A_LWL<436> A_LWL<435> A_LWL<434> A_LWL<433> A_LWL<432> A_LWL<431> A_LWL<430> A_LWL<429> A_LWL<428> A_LWL<427> A_LWL<426> A_LWL<425> A_LWL<424> A_LWL<423> A_LWL<422> A_LWL<421> A_LWL<420> A_LWL<419> A_LWL<418> A_LWL<417> A_LWL<416> A_LWL<415> A_LWL<414> A_LWL<413> A_LWL<412> A_LWL<411> A_LWL<410> A_LWL<409> A_LWL<408> A_LWL<407> A_LWL<406> A_LWL<405> A_LWL<404> A_LWL<403> A_LWL<402> A_LWL<401> A_LWL<400> A_LWL<399> A_LWL<398> A_LWL<397> A_LWL<396> A_LWL<395> A_LWL<394> A_LWL<393> A_LWL<392> A_LWL<391> A_LWL<390> A_LWL<389> A_LWL<388> A_LWL<387> A_LWL<386> A_LWL<385> A_LWL<384> A_LWL<383> A_LWL<382> A_LWL<381> A_LWL<380> A_LWL<379> A_LWL<378> A_LWL<377> A_LWL<376> A_LWL<375> A_LWL<374> A_LWL<373> A_LWL<372> A_LWL<371> A_LWL<370> A_LWL<369> A_LWL<368> A_LWL<367> A_LWL<366> A_LWL<365> A_LWL<364> A_LWL<363> A_LWL<362> A_LWL<361> A_LWL<360> A_LWL<359> A_LWL<358> A_LWL<357> A_LWL<356> A_LWL<355> A_LWL<354> A_LWL<353> A_LWL<352> A_LWL<351> A_LWL<350> A_LWL<349> A_LWL<348> A_LWL<347> A_LWL<346> A_LWL<345> A_LWL<344> A_LWL<343> A_LWL<342> A_LWL<341> A_LWL<340> A_LWL<339> A_LWL<338> A_LWL<337> A_LWL<336> A_LWL<335> A_LWL<334> A_LWL<333> A_LWL<332> A_LWL<331> A_LWL<330> A_LWL<329> A_LWL<328> A_LWL<327> A_LWL<326> A_LWL<325> A_LWL<324> A_LWL<323> A_LWL<322> A_LWL<321> A_LWL<320> A_LWL<319> A_LWL<318> A_LWL<317> A_LWL<316> A_LWL<315> A_LWL<314> A_LWL<313> A_LWL<312> A_LWL<311> A_LWL<310> A_LWL<309> A_LWL<308> A_LWL<307> A_LWL<306> A_LWL<305> A_LWL<304> A_LWL<303> A_LWL<302> A_LWL<301> A_LWL<300> A_LWL<299> A_LWL<298> A_LWL<297> A_LWL<296> A_LWL<295> A_LWL<294> A_LWL<293> A_LWL<292> A_LWL<291> A_LWL<290> A_LWL<289> A_LWL<288> A_LWL<287> A_LWL<286> A_LWL<285> A_LWL<284> A_LWL<283> A_LWL<282> A_LWL<281> A_LWL<280> A_LWL<279> A_LWL<278> A_LWL<277> A_LWL<276> A_LWL<275> A_LWL<274> A_LWL<273> A_LWL<272> A_LWL<271> A_LWL<270> A_LWL<269> A_LWL<268> A_LWL<267> A_LWL<266> A_LWL<265> A_LWL<264> A_LWL<263> A_LWL<262> A_LWL<261> A_LWL<260> A_LWL<259> A_LWL<258> A_LWL<257> A_LWL<256> A_LWL<255> A_LWL<254> A_LWL<253> A_LWL<252> A_LWL<251> A_LWL<250> A_LWL<249> A_LWL<248> A_LWL<247> A_LWL<246> A_LWL<245> A_LWL<244> A_LWL<243> A_LWL<242> A_LWL<241> A_LWL<240> A_LWL<239> A_LWL<238> A_LWL<237> A_LWL<236> A_LWL<235> A_LWL<234> A_LWL<233> A_LWL<232> A_LWL<231> A_LWL<230> A_LWL<229> A_LWL<228> A_LWL<227> A_LWL<226> A_LWL<225> A_LWL<224> A_LWL<223> A_LWL<222> A_LWL<221> A_LWL<220> A_LWL<219> A_LWL<218> A_LWL<217> A_LWL<216> A_LWL<215> A_LWL<214> A_LWL<213> A_LWL<212> A_LWL<211> A_LWL<210> A_LWL<209> A_LWL<208> A_LWL<207> A_LWL<206> A_LWL<205> A_LWL<204> A_LWL<203> A_LWL<202> A_LWL<201> A_LWL<200> A_LWL<199> A_LWL<198> A_LWL<197> A_LWL<196> A_LWL<195> A_LWL<194> A_LWL<193> A_LWL<192> A_LWL<191> A_LWL<190> A_LWL<189> A_LWL<188> A_LWL<187> A_LWL<186> A_LWL<185> A_LWL<184> A_LWL<183> A_LWL<182> A_LWL<181> A_LWL<180> A_LWL<179> A_LWL<178> A_LWL<177> A_LWL<176> A_LWL<175> A_LWL<174> A_LWL<173> A_LWL<172> A_LWL<171> A_LWL<170> A_LWL<169> A_LWL<168> A_LWL<167> A_LWL<166> A_LWL<165> A_LWL<164> A_LWL<163> A_LWL<162> A_LWL<161> A_LWL<160> A_LWL<159> A_LWL<158> A_LWL<157> A_LWL<156> A_LWL<155> A_LWL<154> A_LWL<153> A_LWL<152> A_LWL<151> A_LWL<150> A_LWL<149> A_LWL<148> A_LWL<147> A_LWL<146> A_LWL<145> A_LWL<144> A_LWL<143> A_LWL<142> A_LWL<141> A_LWL<140> A_LWL<139> A_LWL<138> A_LWL<137> A_LWL<136> A_LWL<135> A_LWL<134> A_LWL<133> A_LWL<132> A_LWL<131> A_LWL<130> A_LWL<129> A_LWL<128> A_LWL<127> A_LWL<126> A_LWL<125> A_LWL<124> A_LWL<123> A_LWL<122> A_LWL<121> A_LWL<120> A_LWL<119> A_LWL<118> A_LWL<117> A_LWL<116> A_LWL<115> A_LWL<114> A_LWL<113> A_LWL<112> A_LWL<111> A_LWL<110> A_LWL<109> A_LWL<108> A_LWL<107> A_LWL<106> A_LWL<105> A_LWL<104> A_LWL<103> A_LWL<102> A_LWL<101> A_LWL<100> A_LWL<99> A_LWL<98> A_LWL<97> A_LWL<96> A_LWL<95> A_LWL<94> A_LWL<93> A_LWL<92> A_LWL<91> A_LWL<90> A_LWL<89> A_LWL<88> A_LWL<87> A_LWL<86> A_LWL<85> A_LWL<84> A_LWL<83> A_LWL<82> A_LWL<81> A_LWL<80> A_LWL<79> A_LWL<78> A_LWL<77> A_LWL<76> A_LWL<75> A_LWL<74> A_LWL<73> A_LWL<72> A_LWL<71> A_LWL<70> A_LWL<69> A_LWL<68> A_LWL<67> A_LWL<66> A_LWL<65> A_LWL<64> A_LWL<63> A_LWL<62> A_LWL<61> A_LWL<60> A_LWL<59> A_LWL<58> A_LWL<57> A_LWL<56> A_LWL<55> A_LWL<54> A_LWL<53> A_LWL<52> A_LWL<51> A_LWL<50> A_LWL<49> A_LWL<48> A_LWL<47> A_LWL<46> A_LWL<45> A_LWL<44> A_LWL<43> A_LWL<42> A_LWL<41> A_LWL<40> A_LWL<39> A_LWL<38> A_LWL<37> A_LWL<36> A_LWL<35> A_LWL<34> A_LWL<33> A_LWL<32> A_LWL<31> A_LWL<30> A_LWL<29> A_LWL<28> A_LWL<27> A_LWL<26> A_LWL<25> A_LWL<24> A_LWL<23> A_LWL<22> A_LWL<21> A_LWL<20> A_LWL<19> A_LWL<18> A_LWL<17> A_LWL<16> A_LWL<15> A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<511> A_RWL<510> A_RWL<509> A_RWL<508> A_RWL<507> A_RWL<506> A_RWL<505> A_RWL<504> A_RWL<503> A_RWL<502> A_RWL<501> A_RWL<500> A_RWL<499> A_RWL<498> A_RWL<497> A_RWL<496> A_RWL<495> A_RWL<494> A_RWL<493> A_RWL<492> A_RWL<491> A_RWL<490> A_RWL<489> A_RWL<488> A_RWL<487> A_RWL<486> A_RWL<485> A_RWL<484> A_RWL<483> A_RWL<482> A_RWL<481> A_RWL<480> A_RWL<479> A_RWL<478> A_RWL<477> A_RWL<476> A_RWL<475> A_RWL<474> A_RWL<473> A_RWL<472> A_RWL<471> A_RWL<470> A_RWL<469> A_RWL<468> A_RWL<467> A_RWL<466> A_RWL<465> A_RWL<464> A_RWL<463> A_RWL<462> A_RWL<461> A_RWL<460> A_RWL<459> A_RWL<458> A_RWL<457> A_RWL<456> A_RWL<455> A_RWL<454> A_RWL<453> A_RWL<452> A_RWL<451> A_RWL<450> A_RWL<449> A_RWL<448> A_RWL<447> A_RWL<446> A_RWL<445> A_RWL<444> A_RWL<443> A_RWL<442> A_RWL<441> A_RWL<440> A_RWL<439> A_RWL<438> A_RWL<437> A_RWL<436> A_RWL<435> A_RWL<434> A_RWL<433> A_RWL<432> A_RWL<431> A_RWL<430> A_RWL<429> A_RWL<428> A_RWL<427> A_RWL<426> A_RWL<425> A_RWL<424> A_RWL<423> A_RWL<422> A_RWL<421> A_RWL<420> A_RWL<419> A_RWL<418> A_RWL<417> A_RWL<416> A_RWL<415> A_RWL<414> A_RWL<413> A_RWL<412> A_RWL<411> A_RWL<410> A_RWL<409> A_RWL<408> A_RWL<407> A_RWL<406> A_RWL<405> A_RWL<404> A_RWL<403> A_RWL<402> A_RWL<401> A_RWL<400> A_RWL<399> A_RWL<398> A_RWL<397> A_RWL<396> A_RWL<395> A_RWL<394> A_RWL<393> A_RWL<392> A_RWL<391> A_RWL<390> A_RWL<389> A_RWL<388> A_RWL<387> A_RWL<386> A_RWL<385> A_RWL<384> A_RWL<383> A_RWL<382> A_RWL<381> A_RWL<380> A_RWL<379> A_RWL<378> A_RWL<377> A_RWL<376> A_RWL<375> A_RWL<374> A_RWL<373> A_RWL<372> A_RWL<371> A_RWL<370> A_RWL<369> A_RWL<368> A_RWL<367> A_RWL<366> A_RWL<365> A_RWL<364> A_RWL<363> A_RWL<362> A_RWL<361> A_RWL<360> A_RWL<359> A_RWL<358> A_RWL<357> A_RWL<356> A_RWL<355> A_RWL<354> A_RWL<353> A_RWL<352> A_RWL<351> A_RWL<350> A_RWL<349> A_RWL<348> A_RWL<347> A_RWL<346> A_RWL<345> A_RWL<344> A_RWL<343> A_RWL<342> A_RWL<341> A_RWL<340> A_RWL<339> A_RWL<338> A_RWL<337> A_RWL<336> A_RWL<335> A_RWL<334> A_RWL<333> A_RWL<332> A_RWL<331> A_RWL<330> A_RWL<329> A_RWL<328> A_RWL<327> A_RWL<326> A_RWL<325> A_RWL<324> A_RWL<323> A_RWL<322> A_RWL<321> A_RWL<320> A_RWL<319> A_RWL<318> A_RWL<317> A_RWL<316> A_RWL<315> A_RWL<314> A_RWL<313> A_RWL<312> A_RWL<311> A_RWL<310> A_RWL<309> A_RWL<308> A_RWL<307> A_RWL<306> A_RWL<305> A_RWL<304> A_RWL<303> A_RWL<302> A_RWL<301> A_RWL<300> A_RWL<299> A_RWL<298> A_RWL<297> A_RWL<296> A_RWL<295> A_RWL<294> A_RWL<293> A_RWL<292> A_RWL<291> A_RWL<290> A_RWL<289> A_RWL<288> A_RWL<287> A_RWL<286> A_RWL<285> A_RWL<284> A_RWL<283> A_RWL<282> A_RWL<281> A_RWL<280> A_RWL<279> A_RWL<278> A_RWL<277> A_RWL<276> A_RWL<275> A_RWL<274> A_RWL<273> A_RWL<272> A_RWL<271> A_RWL<270> A_RWL<269> A_RWL<268> A_RWL<267> A_RWL<266> A_RWL<265> A_RWL<264> A_RWL<263> A_RWL<262> A_RWL<261> A_RWL<260> A_RWL<259> A_RWL<258> A_RWL<257> A_RWL<256> A_RWL<255> A_RWL<254> A_RWL<253> A_RWL<252> A_RWL<251> A_RWL<250> A_RWL<249> A_RWL<248> A_RWL<247> A_RWL<246> A_RWL<245> A_RWL<244> A_RWL<243> A_RWL<242> A_RWL<241> A_RWL<240> A_RWL<239> A_RWL<238> A_RWL<237> A_RWL<236> A_RWL<235> A_RWL<234> A_RWL<233> A_RWL<232> A_RWL<231> A_RWL<230> A_RWL<229> A_RWL<228> A_RWL<227> A_RWL<226> A_RWL<225> A_RWL<224> A_RWL<223> A_RWL<222> A_RWL<221> A_RWL<220> A_RWL<219> A_RWL<218> A_RWL<217> A_RWL<216> A_RWL<215> A_RWL<214> A_RWL<213> A_RWL<212> A_RWL<211> A_RWL<210> A_RWL<209> A_RWL<208> A_RWL<207> A_RWL<206> A_RWL<205> A_RWL<204> A_RWL<203> A_RWL<202> A_RWL<201> A_RWL<200> A_RWL<199> A_RWL<198> A_RWL<197> A_RWL<196> A_RWL<195> A_RWL<194> A_RWL<193> A_RWL<192> A_RWL<191> A_RWL<190> A_RWL<189> A_RWL<188> A_RWL<187> A_RWL<186> A_RWL<185> A_RWL<184> A_RWL<183> A_RWL<182> A_RWL<181> A_RWL<180> A_RWL<179> A_RWL<178> A_RWL<177> A_RWL<176> A_RWL<175> A_RWL<174> A_RWL<173> A_RWL<172> A_RWL<171> A_RWL<170> A_RWL<169> A_RWL<168> A_RWL<167> A_RWL<166> A_RWL<165> A_RWL<164> A_RWL<163> A_RWL<162> A_RWL<161> A_RWL<160> A_RWL<159> A_RWL<158> A_RWL<157> A_RWL<156> A_RWL<155> A_RWL<154> A_RWL<153> A_RWL<152> A_RWL<151> A_RWL<150> A_RWL<149> A_RWL<148> A_RWL<147> A_RWL<146> A_RWL<145> A_RWL<144> A_RWL<143> A_RWL<142> A_RWL<141> A_RWL<140> A_RWL<139> A_RWL<138> A_RWL<137> A_RWL<136> A_RWL<135> A_RWL<134> A_RWL<133> A_RWL<132> A_RWL<131> A_RWL<130> A_RWL<129> A_RWL<128> A_RWL<127> A_RWL<126> A_RWL<125> A_RWL<124> A_RWL<123> A_RWL<122> A_RWL<121> A_RWL<120> A_RWL<119> A_RWL<118> A_RWL<117> A_RWL<116> A_RWL<115> A_RWL<114> A_RWL<113> A_RWL<112> A_RWL<111> A_RWL<110> A_RWL<109> A_RWL<108> A_RWL<107> A_RWL<106> A_RWL<105> A_RWL<104> A_RWL<103> A_RWL<102> A_RWL<101> A_RWL<100> A_RWL<99> A_RWL<98> A_RWL<97> A_RWL<96> A_RWL<95> A_RWL<94> A_RWL<93> A_RWL<92> A_RWL<91> A_RWL<90> A_RWL<89> A_RWL<88> A_RWL<87> A_RWL<86> A_RWL<85> A_RWL<84> A_RWL<83> A_RWL<82> A_RWL<81> A_RWL<80> A_RWL<79> A_RWL<78> A_RWL<77> A_RWL<76> A_RWL<75> A_RWL<74> A_RWL<73> A_RWL<72> A_RWL<71> A_RWL<70> A_RWL<69> A_RWL<68> A_RWL<67> A_RWL<66> A_RWL<65> A_RWL<64> A_RWL<63> A_RWL<62> A_RWL<61> A_RWL<60> A_RWL<59> A_RWL<58> A_RWL<57> A_RWL<56> A_RWL<55> A_RWL<54> A_RWL<53> A_RWL<52> A_RWL<51> A_RWL<50> A_RWL<49> A_RWL<48> A_RWL<47> A_RWL<46> A_RWL<45> A_RWL<44> A_RWL<43> A_RWL<42> A_RWL<41> A_RWL<40> A_RWL<39> A_RWL<38> A_RWL<37> A_RWL<36> A_RWL<35> A_RWL<34> A_RWL<33> A_RWL<32> A_RWL<31> A_RWL<30> A_RWL<29> A_RWL<28> A_RWL<27> A_RWL<26> A_RWL<25> A_RWL<24> A_RWL<23> A_RWL<22> A_RWL<21> A_RWL<20> A_RWL<19> A_RWL<18> A_RWL<17> A_RWL<16> A_RWL<15> A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE VSS
XRAM<32> A_BLC<61> A_BLC<60> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT<61> A_BLT<60> A_BLT_TOP<1> A_BLT_TOP<0> A_LWL<511> A_LWL<510> A_LWL<509> A_LWL<508> A_LWL<507> A_LWL<506> A_LWL<505> A_LWL<504> A_LWL<503> A_LWL<502> A_LWL<501> A_LWL<500> A_LWL<499> A_LWL<498> A_LWL<497> A_LWL<496> A_RWL<511> A_RWL<510> A_RWL<509> A_RWL<508> A_RWL<507> A_RWL<506> A_RWL<505> A_RWL<504> A_RWL<503> A_RWL<502> A_RWL<501> A_RWL<500> A_RWL<499> A_RWL<498> A_RWL<497> A_RWL<496> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<31> A_BLC<59> A_BLC<58> A_BLC<61> A_BLC<60> A_BLT<59> A_BLT<58> A_BLT<61> A_BLT<60> A_LWL<495> A_LWL<494> A_LWL<493> A_LWL<492> A_LWL<491> A_LWL<490> A_LWL<489> A_LWL<488> A_LWL<487> A_LWL<486> A_LWL<485> A_LWL<484> A_LWL<483> A_LWL<482> A_LWL<481> A_LWL<480> A_RWL<495> A_RWL<494> A_RWL<493> A_RWL<492> A_RWL<491> A_RWL<490> A_RWL<489> A_RWL<488> A_RWL<487> A_RWL<486> A_RWL<485> A_RWL<484> A_RWL<483> A_RWL<482> A_RWL<481> A_RWL<480> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<30> A_BLC<57> A_BLC<56> A_BLC<59> A_BLC<58> A_BLT<57> A_BLT<56> A_BLT<59> A_BLT<58> A_LWL<479> A_LWL<478> A_LWL<477> A_LWL<476> A_LWL<475> A_LWL<474> A_LWL<473> A_LWL<472> A_LWL<471> A_LWL<470> A_LWL<469> A_LWL<468> A_LWL<467> A_LWL<466> A_LWL<465> A_LWL<464> A_RWL<479> A_RWL<478> A_RWL<477> A_RWL<476> A_RWL<475> A_RWL<474> A_RWL<473> A_RWL<472> A_RWL<471> A_RWL<470> A_RWL<469> A_RWL<468> A_RWL<467> A_RWL<466> A_RWL<465> A_RWL<464> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<29> A_BLC<55> A_BLC<54> A_BLC<57> A_BLC<56> A_BLT<55> A_BLT<54> A_BLT<57> A_BLT<56> A_LWL<463> A_LWL<462> A_LWL<461> A_LWL<460> A_LWL<459> A_LWL<458> A_LWL<457> A_LWL<456> A_LWL<455> A_LWL<454> A_LWL<453> A_LWL<452> A_LWL<451> A_LWL<450> A_LWL<449> A_LWL<448> A_RWL<463> A_RWL<462> A_RWL<461> A_RWL<460> A_RWL<459> A_RWL<458> A_RWL<457> A_RWL<456> A_RWL<455> A_RWL<454> A_RWL<453> A_RWL<452> A_RWL<451> A_RWL<450> A_RWL<449> A_RWL<448> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<28> A_BLC<53> A_BLC<52> A_BLC<55> A_BLC<54> A_BLT<53> A_BLT<52> A_BLT<55> A_BLT<54> A_LWL<447> A_LWL<446> A_LWL<445> A_LWL<444> A_LWL<443> A_LWL<442> A_LWL<441> A_LWL<440> A_LWL<439> A_LWL<438> A_LWL<437> A_LWL<436> A_LWL<435> A_LWL<434> A_LWL<433> A_LWL<432> A_RWL<447> A_RWL<446> A_RWL<445> A_RWL<444> A_RWL<443> A_RWL<442> A_RWL<441> A_RWL<440> A_RWL<439> A_RWL<438> A_RWL<437> A_RWL<436> A_RWL<435> A_RWL<434> A_RWL<433> A_RWL<432> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<27> A_BLC<51> A_BLC<50> A_BLC<53> A_BLC<52> A_BLT<51> A_BLT<50> A_BLT<53> A_BLT<52> A_LWL<431> A_LWL<430> A_LWL<429> A_LWL<428> A_LWL<427> A_LWL<426> A_LWL<425> A_LWL<424> A_LWL<423> A_LWL<422> A_LWL<421> A_LWL<420> A_LWL<419> A_LWL<418> A_LWL<417> A_LWL<416> A_RWL<431> A_RWL<430> A_RWL<429> A_RWL<428> A_RWL<427> A_RWL<426> A_RWL<425> A_RWL<424> A_RWL<423> A_RWL<422> A_RWL<421> A_RWL<420> A_RWL<419> A_RWL<418> A_RWL<417> A_RWL<416> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<26> A_BLC<49> A_BLC<48> A_BLC<51> A_BLC<50> A_BLT<49> A_BLT<48> A_BLT<51> A_BLT<50> A_LWL<415> A_LWL<414> A_LWL<413> A_LWL<412> A_LWL<411> A_LWL<410> A_LWL<409> A_LWL<408> A_LWL<407> A_LWL<406> A_LWL<405> A_LWL<404> A_LWL<403> A_LWL<402> A_LWL<401> A_LWL<400> A_RWL<415> A_RWL<414> A_RWL<413> A_RWL<412> A_RWL<411> A_RWL<410> A_RWL<409> A_RWL<408> A_RWL<407> A_RWL<406> A_RWL<405> A_RWL<404> A_RWL<403> A_RWL<402> A_RWL<401> A_RWL<400> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<25> A_BLC<47> A_BLC<46> A_BLC<49> A_BLC<48> A_BLT<47> A_BLT<46> A_BLT<49> A_BLT<48> A_LWL<399> A_LWL<398> A_LWL<397> A_LWL<396> A_LWL<395> A_LWL<394> A_LWL<393> A_LWL<392> A_LWL<391> A_LWL<390> A_LWL<389> A_LWL<388> A_LWL<387> A_LWL<386> A_LWL<385> A_LWL<384> A_RWL<399> A_RWL<398> A_RWL<397> A_RWL<396> A_RWL<395> A_RWL<394> A_RWL<393> A_RWL<392> A_RWL<391> A_RWL<390> A_RWL<389> A_RWL<388> A_RWL<387> A_RWL<386> A_RWL<385> A_RWL<384> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<24> A_BLC<45> A_BLC<44> A_BLC<47> A_BLC<46> A_BLT<45> A_BLT<44> A_BLT<47> A_BLT<46> A_LWL<383> A_LWL<382> A_LWL<381> A_LWL<380> A_LWL<379> A_LWL<378> A_LWL<377> A_LWL<376> A_LWL<375> A_LWL<374> A_LWL<373> A_LWL<372> A_LWL<371> A_LWL<370> A_LWL<369> A_LWL<368> A_RWL<383> A_RWL<382> A_RWL<381> A_RWL<380> A_RWL<379> A_RWL<378> A_RWL<377> A_RWL<376> A_RWL<375> A_RWL<374> A_RWL<373> A_RWL<372> A_RWL<371> A_RWL<370> A_RWL<369> A_RWL<368> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<23> A_BLC<43> A_BLC<42> A_BLC<45> A_BLC<44> A_BLT<43> A_BLT<42> A_BLT<45> A_BLT<44> A_LWL<367> A_LWL<366> A_LWL<365> A_LWL<364> A_LWL<363> A_LWL<362> A_LWL<361> A_LWL<360> A_LWL<359> A_LWL<358> A_LWL<357> A_LWL<356> A_LWL<355> A_LWL<354> A_LWL<353> A_LWL<352> A_RWL<367> A_RWL<366> A_RWL<365> A_RWL<364> A_RWL<363> A_RWL<362> A_RWL<361> A_RWL<360> A_RWL<359> A_RWL<358> A_RWL<357> A_RWL<356> A_RWL<355> A_RWL<354> A_RWL<353> A_RWL<352> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<22> A_BLC<41> A_BLC<40> A_BLC<43> A_BLC<42> A_BLT<41> A_BLT<40> A_BLT<43> A_BLT<42> A_LWL<351> A_LWL<350> A_LWL<349> A_LWL<348> A_LWL<347> A_LWL<346> A_LWL<345> A_LWL<344> A_LWL<343> A_LWL<342> A_LWL<341> A_LWL<340> A_LWL<339> A_LWL<338> A_LWL<337> A_LWL<336> A_RWL<351> A_RWL<350> A_RWL<349> A_RWL<348> A_RWL<347> A_RWL<346> A_RWL<345> A_RWL<344> A_RWL<343> A_RWL<342> A_RWL<341> A_RWL<340> A_RWL<339> A_RWL<338> A_RWL<337> A_RWL<336> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<21> A_BLC<39> A_BLC<38> A_BLC<41> A_BLC<40> A_BLT<39> A_BLT<38> A_BLT<41> A_BLT<40> A_LWL<335> A_LWL<334> A_LWL<333> A_LWL<332> A_LWL<331> A_LWL<330> A_LWL<329> A_LWL<328> A_LWL<327> A_LWL<326> A_LWL<325> A_LWL<324> A_LWL<323> A_LWL<322> A_LWL<321> A_LWL<320> A_RWL<335> A_RWL<334> A_RWL<333> A_RWL<332> A_RWL<331> A_RWL<330> A_RWL<329> A_RWL<328> A_RWL<327> A_RWL<326> A_RWL<325> A_RWL<324> A_RWL<323> A_RWL<322> A_RWL<321> A_RWL<320> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<20> A_BLC<37> A_BLC<36> A_BLC<39> A_BLC<38> A_BLT<37> A_BLT<36> A_BLT<39> A_BLT<38> A_LWL<319> A_LWL<318> A_LWL<317> A_LWL<316> A_LWL<315> A_LWL<314> A_LWL<313> A_LWL<312> A_LWL<311> A_LWL<310> A_LWL<309> A_LWL<308> A_LWL<307> A_LWL<306> A_LWL<305> A_LWL<304> A_RWL<319> A_RWL<318> A_RWL<317> A_RWL<316> A_RWL<315> A_RWL<314> A_RWL<313> A_RWL<312> A_RWL<311> A_RWL<310> A_RWL<309> A_RWL<308> A_RWL<307> A_RWL<306> A_RWL<305> A_RWL<304> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<19> A_BLC<35> A_BLC<34> A_BLC<37> A_BLC<36> A_BLT<35> A_BLT<34> A_BLT<37> A_BLT<36> A_LWL<303> A_LWL<302> A_LWL<301> A_LWL<300> A_LWL<299> A_LWL<298> A_LWL<297> A_LWL<296> A_LWL<295> A_LWL<294> A_LWL<293> A_LWL<292> A_LWL<291> A_LWL<290> A_LWL<289> A_LWL<288> A_RWL<303> A_RWL<302> A_RWL<301> A_RWL<300> A_RWL<299> A_RWL<298> A_RWL<297> A_RWL<296> A_RWL<295> A_RWL<294> A_RWL<293> A_RWL<292> A_RWL<291> A_RWL<290> A_RWL<289> A_RWL<288> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<18> A_BLC<33> A_BLC<32> A_BLC<35> A_BLC<34> A_BLT<33> A_BLT<32> A_BLT<35> A_BLT<34> A_LWL<287> A_LWL<286> A_LWL<285> A_LWL<284> A_LWL<283> A_LWL<282> A_LWL<281> A_LWL<280> A_LWL<279> A_LWL<278> A_LWL<277> A_LWL<276> A_LWL<275> A_LWL<274> A_LWL<273> A_LWL<272> A_RWL<287> A_RWL<286> A_RWL<285> A_RWL<284> A_RWL<283> A_RWL<282> A_RWL<281> A_RWL<280> A_RWL<279> A_RWL<278> A_RWL<277> A_RWL<276> A_RWL<275> A_RWL<274> A_RWL<273> A_RWL<272> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<17> A_BLC<31> A_BLC<30> A_BLC<33> A_BLC<32> A_BLT<31> A_BLT<30> A_BLT<33> A_BLT<32> A_LWL<271> A_LWL<270> A_LWL<269> A_LWL<268> A_LWL<267> A_LWL<266> A_LWL<265> A_LWL<264> A_LWL<263> A_LWL<262> A_LWL<261> A_LWL<260> A_LWL<259> A_LWL<258> A_LWL<257> A_LWL<256> A_RWL<271> A_RWL<270> A_RWL<269> A_RWL<268> A_RWL<267> A_RWL<266> A_RWL<265> A_RWL<264> A_RWL<263> A_RWL<262> A_RWL<261> A_RWL<260> A_RWL<259> A_RWL<258> A_RWL<257> A_RWL<256> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<16> A_BLC<29> A_BLC<28> A_BLC<31> A_BLC<30> A_BLT<29> A_BLT<28> A_BLT<31> A_BLT<30> A_LWL<255> A_LWL<254> A_LWL<253> A_LWL<252> A_LWL<251> A_LWL<250> A_LWL<249> A_LWL<248> A_LWL<247> A_LWL<246> A_LWL<245> A_LWL<244> A_LWL<243> A_LWL<242> A_LWL<241> A_LWL<240> A_RWL<255> A_RWL<254> A_RWL<253> A_RWL<252> A_RWL<251> A_RWL<250> A_RWL<249> A_RWL<248> A_RWL<247> A_RWL<246> A_RWL<245> A_RWL<244> A_RWL<243> A_RWL<242> A_RWL<241> A_RWL<240> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<15> A_BLC<27> A_BLC<26> A_BLC<29> A_BLC<28> A_BLT<27> A_BLT<26> A_BLT<29> A_BLT<28> A_LWL<239> A_LWL<238> A_LWL<237> A_LWL<236> A_LWL<235> A_LWL<234> A_LWL<233> A_LWL<232> A_LWL<231> A_LWL<230> A_LWL<229> A_LWL<228> A_LWL<227> A_LWL<226> A_LWL<225> A_LWL<224> A_RWL<239> A_RWL<238> A_RWL<237> A_RWL<236> A_RWL<235> A_RWL<234> A_RWL<233> A_RWL<232> A_RWL<231> A_RWL<230> A_RWL<229> A_RWL<228> A_RWL<227> A_RWL<226> A_RWL<225> A_RWL<224> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<14> A_BLC<25> A_BLC<24> A_BLC<27> A_BLC<26> A_BLT<25> A_BLT<24> A_BLT<27> A_BLT<26> A_LWL<223> A_LWL<222> A_LWL<221> A_LWL<220> A_LWL<219> A_LWL<218> A_LWL<217> A_LWL<216> A_LWL<215> A_LWL<214> A_LWL<213> A_LWL<212> A_LWL<211> A_LWL<210> A_LWL<209> A_LWL<208> A_RWL<223> A_RWL<222> A_RWL<221> A_RWL<220> A_RWL<219> A_RWL<218> A_RWL<217> A_RWL<216> A_RWL<215> A_RWL<214> A_RWL<213> A_RWL<212> A_RWL<211> A_RWL<210> A_RWL<209> A_RWL<208> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<13> A_BLC<23> A_BLC<22> A_BLC<25> A_BLC<24> A_BLT<23> A_BLT<22> A_BLT<25> A_BLT<24> A_LWL<207> A_LWL<206> A_LWL<205> A_LWL<204> A_LWL<203> A_LWL<202> A_LWL<201> A_LWL<200> A_LWL<199> A_LWL<198> A_LWL<197> A_LWL<196> A_LWL<195> A_LWL<194> A_LWL<193> A_LWL<192> A_RWL<207> A_RWL<206> A_RWL<205> A_RWL<204> A_RWL<203> A_RWL<202> A_RWL<201> A_RWL<200> A_RWL<199> A_RWL<198> A_RWL<197> A_RWL<196> A_RWL<195> A_RWL<194> A_RWL<193> A_RWL<192> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<12> A_BLC<21> A_BLC<20> A_BLC<23> A_BLC<22> A_BLT<21> A_BLT<20> A_BLT<23> A_BLT<22> A_LWL<191> A_LWL<190> A_LWL<189> A_LWL<188> A_LWL<187> A_LWL<186> A_LWL<185> A_LWL<184> A_LWL<183> A_LWL<182> A_LWL<181> A_LWL<180> A_LWL<179> A_LWL<178> A_LWL<177> A_LWL<176> A_RWL<191> A_RWL<190> A_RWL<189> A_RWL<188> A_RWL<187> A_RWL<186> A_RWL<185> A_RWL<184> A_RWL<183> A_RWL<182> A_RWL<181> A_RWL<180> A_RWL<179> A_RWL<178> A_RWL<177> A_RWL<176> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<11> A_BLC<19> A_BLC<18> A_BLC<21> A_BLC<20> A_BLT<19> A_BLT<18> A_BLT<21> A_BLT<20> A_LWL<175> A_LWL<174> A_LWL<173> A_LWL<172> A_LWL<171> A_LWL<170> A_LWL<169> A_LWL<168> A_LWL<167> A_LWL<166> A_LWL<165> A_LWL<164> A_LWL<163> A_LWL<162> A_LWL<161> A_LWL<160> A_RWL<175> A_RWL<174> A_RWL<173> A_RWL<172> A_RWL<171> A_RWL<170> A_RWL<169> A_RWL<168> A_RWL<167> A_RWL<166> A_RWL<165> A_RWL<164> A_RWL<163> A_RWL<162> A_RWL<161> A_RWL<160> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<10> A_BLC<17> A_BLC<16> A_BLC<19> A_BLC<18> A_BLT<17> A_BLT<16> A_BLT<19> A_BLT<18> A_LWL<159> A_LWL<158> A_LWL<157> A_LWL<156> A_LWL<155> A_LWL<154> A_LWL<153> A_LWL<152> A_LWL<151> A_LWL<150> A_LWL<149> A_LWL<148> A_LWL<147> A_LWL<146> A_LWL<145> A_LWL<144> A_RWL<159> A_RWL<158> A_RWL<157> A_RWL<156> A_RWL<155> A_RWL<154> A_RWL<153> A_RWL<152> A_RWL<151> A_RWL<150> A_RWL<149> A_RWL<148> A_RWL<147> A_RWL<146> A_RWL<145> A_RWL<144> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<9> A_BLC<15> A_BLC<14> A_BLC<17> A_BLC<16> A_BLT<15> A_BLT<14> A_BLT<17> A_BLT<16> A_LWL<143> A_LWL<142> A_LWL<141> A_LWL<140> A_LWL<139> A_LWL<138> A_LWL<137> A_LWL<136> A_LWL<135> A_LWL<134> A_LWL<133> A_LWL<132> A_LWL<131> A_LWL<130> A_LWL<129> A_LWL<128> A_RWL<143> A_RWL<142> A_RWL<141> A_RWL<140> A_RWL<139> A_RWL<138> A_RWL<137> A_RWL<136> A_RWL<135> A_RWL<134> A_RWL<133> A_RWL<132> A_RWL<131> A_RWL<130> A_RWL<129> A_RWL<128> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<8> A_BLC<13> A_BLC<12> A_BLC<15> A_BLC<14> A_BLT<13> A_BLT<12> A_BLT<15> A_BLT<14> A_LWL<127> A_LWL<126> A_LWL<125> A_LWL<124> A_LWL<123> A_LWL<122> A_LWL<121> A_LWL<120> A_LWL<119> A_LWL<118> A_LWL<117> A_LWL<116> A_LWL<115> A_LWL<114> A_LWL<113> A_LWL<112> A_RWL<127> A_RWL<126> A_RWL<125> A_RWL<124> A_RWL<123> A_RWL<122> A_RWL<121> A_RWL<120> A_RWL<119> A_RWL<118> A_RWL<117> A_RWL<116> A_RWL<115> A_RWL<114> A_RWL<113> A_RWL<112> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<7> A_BLC<11> A_BLC<10> A_BLC<13> A_BLC<12> A_BLT<11> A_BLT<10> A_BLT<13> A_BLT<12> A_LWL<111> A_LWL<110> A_LWL<109> A_LWL<108> A_LWL<107> A_LWL<106> A_LWL<105> A_LWL<104> A_LWL<103> A_LWL<102> A_LWL<101> A_LWL<100> A_LWL<99> A_LWL<98> A_LWL<97> A_LWL<96> A_RWL<111> A_RWL<110> A_RWL<109> A_RWL<108> A_RWL<107> A_RWL<106> A_RWL<105> A_RWL<104> A_RWL<103> A_RWL<102> A_RWL<101> A_RWL<100> A_RWL<99> A_RWL<98> A_RWL<97> A_RWL<96> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<6> A_BLC<9> A_BLC<8> A_BLC<11> A_BLC<10> A_BLT<9> A_BLT<8> A_BLT<11> A_BLT<10> A_LWL<95> A_LWL<94> A_LWL<93> A_LWL<92> A_LWL<91> A_LWL<90> A_LWL<89> A_LWL<88> A_LWL<87> A_LWL<86> A_LWL<85> A_LWL<84> A_LWL<83> A_LWL<82> A_LWL<81> A_LWL<80> A_RWL<95> A_RWL<94> A_RWL<93> A_RWL<92> A_RWL<91> A_RWL<90> A_RWL<89> A_RWL<88> A_RWL<87> A_RWL<86> A_RWL<85> A_RWL<84> A_RWL<83> A_RWL<82> A_RWL<81> A_RWL<80> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<5> A_BLC<7> A_BLC<6> A_BLC<9> A_BLC<8> A_BLT<7> A_BLT<6> A_BLT<9> A_BLT<8> A_LWL<79> A_LWL<78> A_LWL<77> A_LWL<76> A_LWL<75> A_LWL<74> A_LWL<73> A_LWL<72> A_LWL<71> A_LWL<70> A_LWL<69> A_LWL<68> A_LWL<67> A_LWL<66> A_LWL<65> A_LWL<64> A_RWL<79> A_RWL<78> A_RWL<77> A_RWL<76> A_RWL<75> A_RWL<74> A_RWL<73> A_RWL<72> A_RWL<71> A_RWL<70> A_RWL<69> A_RWL<68> A_RWL<67> A_RWL<66> A_RWL<65> A_RWL<64> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<4> A_BLC<5> A_BLC<4> A_BLC<7> A_BLC<6> A_BLT<5> A_BLT<4> A_BLT<7> A_BLT<6> A_LWL<63> A_LWL<62> A_LWL<61> A_LWL<60> A_LWL<59> A_LWL<58> A_LWL<57> A_LWL<56> A_LWL<55> A_LWL<54> A_LWL<53> A_LWL<52> A_LWL<51> A_LWL<50> A_LWL<49> A_LWL<48> A_RWL<63> A_RWL<62> A_RWL<61> A_RWL<60> A_RWL<59> A_RWL<58> A_RWL<57> A_RWL<56> A_RWL<55> A_RWL<54> A_RWL<53> A_RWL<52> A_RWL<51> A_RWL<50> A_RWL<49> A_RWL<48> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<3> A_BLC<3> A_BLC<2> A_BLC<5> A_BLC<4> A_BLT<3> A_BLT<2> A_BLT<5> A_BLT<4> A_LWL<47> A_LWL<46> A_LWL<45> A_LWL<44> A_LWL<43> A_LWL<42> A_LWL<41> A_LWL<40> A_LWL<39> A_LWL<38> A_LWL<37> A_LWL<36> A_LWL<35> A_LWL<34> A_LWL<33> A_LWL<32> A_RWL<47> A_RWL<46> A_RWL<45> A_RWL<44> A_RWL<43> A_RWL<42> A_RWL<41> A_RWL<40> A_RWL<39> A_RWL<38> A_RWL<37> A_RWL<36> A_RWL<35> A_RWL<34> A_RWL<33> A_RWL<32> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<2> A_BLC<1> A_BLC<0> A_BLC<3> A_BLC<2> A_BLT<1> A_BLT<0> A_BLT<3> A_BLT<2> A_LWL<31> A_LWL<30> A_LWL<29> A_LWL<28> A_LWL<27> A_LWL<26> A_LWL<25> A_LWL<24> A_LWL<23> A_LWL<22> A_LWL<21> A_LWL<20> A_LWL<19> A_LWL<18> A_LWL<17> A_LWL<16> A_RWL<31> A_RWL<30> A_RWL<29> A_RWL<28> A_RWL<27> A_RWL<26> A_RWL<25> A_RWL<24> A_RWL<23> A_RWL<22> A_RWL<21> A_RWL<20> A_RWL<19> A_RWL<18> A_RWL<17> A_RWL<16> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XRAM<1> A_BLC_BOT<1> A_BLC_BOT<0> A_BLC<1> A_BLC<0> A_BLT_BOT<1> A_BLT_BOT<0> A_BLT<1> A_BLT<0> A_LWL<15> A_LWL<14> A_LWL<13> A_LWL<12> A_LWL<11> A_LWL<10> A_LWL<9> A_LWL<8> A_LWL<7> A_LWL<6> A_LWL<5> A_LWL<4> A_LWL<3> A_LWL<2> A_LWL<1> A_LWL<0> A_RWL<15> A_RWL<14> A_RWL<13> A_RWL<12> A_RWL<11> A_RWL<10> A_RWL<9> A_RWL<8> A_RWL<7> A_RWL<6> A_RWL<5> A_RWL<4> A_RWL<3> A_RWL<2> A_RWL<1> A_RWL<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_SRAM
XEDGE<1> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT_TOP<1> A_BLT_TOP<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_TB
XEDGE<0> A_BLC_BOT<1> A_BLC_BOT<0> A_BLT_BOT<1> A_BLT_BOT<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_TB
.ENDS




.SUBCKT RM_IHPSG13_2048x64_c2_1P_MATRIX_pcell_1 A_BLC<127> A_BLC<126> A_BLC<125> A_BLC<124> A_BLC<123> A_BLC<122> A_BLC<121> A_BLC<120> A_BLC<119> A_BLC<118> A_BLC<117> A_BLC<116> A_BLC<115> A_BLC<114> A_BLC<113> A_BLC<112> A_BLC<111> A_BLC<110> A_BLC<109> A_BLC<108> A_BLC<107> A_BLC<106> A_BLC<105> A_BLC<104> A_BLC<103> A_BLC<102> A_BLC<101> A_BLC<100> A_BLC<99> A_BLC<98> A_BLC<97> A_BLC<96> A_BLC<95> A_BLC<94> A_BLC<93> A_BLC<92> A_BLC<91> A_BLC<90> A_BLC<89> A_BLC<88> A_BLC<87> A_BLC<86> A_BLC<85> A_BLC<84> A_BLC<83> A_BLC<82> A_BLC<81> A_BLC<80> A_BLC<79> A_BLC<78> A_BLC<77> A_BLC<76> A_BLC<75> A_BLC<74> A_BLC<73> A_BLC<72> A_BLC<71> A_BLC<70> A_BLC<69> A_BLC<68> A_BLC<67> A_BLC<66> A_BLC<65> A_BLC<64> A_BLC<63> A_BLC<62> A_BLC<61> A_BLC<60> A_BLC<59> A_BLC<58> A_BLC<57> A_BLC<56> A_BLC<55> A_BLC<54> A_BLC<53> A_BLC<52> A_BLC<51> A_BLC<50> A_BLC<49> A_BLC<48> A_BLC<47> A_BLC<46> A_BLC<45> A_BLC<44> A_BLC<43> A_BLC<42> A_BLC<41> A_BLC<40> A_BLC<39> A_BLC<38> A_BLC<37> A_BLC<36> A_BLC<35> A_BLC<34> A_BLC<33> A_BLC<32> A_BLC<31> A_BLC<30> A_BLC<29> A_BLC<28> A_BLC<27> A_BLC<26> A_BLC<25> A_BLC<24> A_BLC<23> A_BLC<22> A_BLC<21> A_BLC<20> A_BLC<19> A_BLC<18> A_BLC<17> A_BLC<16> A_BLC<15> A_BLC<14> A_BLC<13> A_BLC<12> A_BLC<11> A_BLC<10> A_BLC<9> A_BLC<8> A_BLC<7> A_BLC<6> A_BLC<5> A_BLC<4> A_BLC<3> A_BLC<2> A_BLC<1> A_BLC<0> A_BLT<127> A_BLT<126> A_BLT<125> A_BLT<124> A_BLT<123> A_BLT<122> A_BLT<121> A_BLT<120> A_BLT<119> A_BLT<118> A_BLT<117> A_BLT<116> A_BLT<115> A_BLT<114> A_BLT<113> A_BLT<112> A_BLT<111> A_BLT<110> A_BLT<109> A_BLT<108> A_BLT<107> A_BLT<106> A_BLT<105> A_BLT<104> A_BLT<103> A_BLT<102> A_BLT<101> A_BLT<100> A_BLT<99> A_BLT<98> A_BLT<97> A_BLT<96> A_BLT<95> A_BLT<94> A_BLT<93> A_BLT<92> A_BLT<91> A_BLT<90> A_BLT<89> A_BLT<88> A_BLT<87> A_BLT<86> A_BLT<85> A_BLT<84> A_BLT<83> A_BLT<82> A_BLT<81> A_BLT<80> A_BLT<79> A_BLT<78> A_BLT<77> A_BLT<76> A_BLT<75> A_BLT<74> A_BLT<73> A_BLT<72> A_BLT<71> A_BLT<70> A_BLT<69> A_BLT<68> A_BLT<67> A_BLT<66> A_BLT<65> A_BLT<64> A_BLT<63> A_BLT<62> A_BLT<61> A_BLT<60> A_BLT<59> A_BLT<58> A_BLT<57> A_BLT<56> A_BLT<55> A_BLT<54> A_BLT<53> A_BLT<52> A_BLT<51> A_BLT<50> A_BLT<49> A_BLT<48> A_BLT<47> A_BLT<46> A_BLT<45> A_BLT<44> A_BLT<43> A_BLT<42> A_BLT<41> A_BLT<40> A_BLT<39> A_BLT<38> A_BLT<37> A_BLT<36> A_BLT<35> A_BLT<34> A_BLT<33> A_BLT<32> A_BLT<31> A_BLT<30> A_BLT<29> A_BLT<28> A_BLT<27> A_BLT<26> A_BLT<25> A_BLT<24> A_BLT<23> A_BLT<22> A_BLT<21> A_BLT<20> A_BLT<19> A_BLT<18> A_BLT<17> A_BLT<16> A_BLT<15> A_BLT<14> A_BLT<13> A_BLT<12> A_BLT<11> A_BLT<10> A_BLT<9> A_BLT<8> A_BLT<7> A_BLT<6> A_BLT<5> A_BLT<4> A_BLT<3> A_BLT<2> A_BLT<1> A_BLT<0> A_WL<511> A_WL<510> A_WL<509> A_WL<508> A_WL<507> A_WL<506> A_WL<505> A_WL<504> A_WL<503> A_WL<502> A_WL<501> A_WL<500> A_WL<499> A_WL<498> A_WL<497> A_WL<496> A_WL<495> A_WL<494> A_WL<493> A_WL<492> A_WL<491> A_WL<490> A_WL<489> A_WL<488> A_WL<487> A_WL<486> A_WL<485> A_WL<484> A_WL<483> A_WL<482> A_WL<481> A_WL<480> A_WL<479> A_WL<478> A_WL<477> A_WL<476> A_WL<475> A_WL<474> A_WL<473> A_WL<472> A_WL<471> A_WL<470> A_WL<469> A_WL<468> A_WL<467> A_WL<466> A_WL<465> A_WL<464> A_WL<463> A_WL<462> A_WL<461> A_WL<460> A_WL<459> A_WL<458> A_WL<457> A_WL<456> A_WL<455> A_WL<454> A_WL<453> A_WL<452> A_WL<451> A_WL<450> A_WL<449> A_WL<448> A_WL<447> A_WL<446> A_WL<445> A_WL<444> A_WL<443> A_WL<442> A_WL<441> A_WL<440> A_WL<439> A_WL<438> A_WL<437> A_WL<436> A_WL<435> A_WL<434> A_WL<433> A_WL<432> A_WL<431> A_WL<430> A_WL<429> A_WL<428> A_WL<427> A_WL<426> A_WL<425> A_WL<424> A_WL<423> A_WL<422> A_WL<421> A_WL<420> A_WL<419> A_WL<418> A_WL<417> A_WL<416> A_WL<415> A_WL<414> A_WL<413> A_WL<412> A_WL<411> A_WL<410> A_WL<409> A_WL<408> A_WL<407> A_WL<406> A_WL<405> A_WL<404> A_WL<403> A_WL<402> A_WL<401> A_WL<400> A_WL<399> A_WL<398> A_WL<397> A_WL<396> A_WL<395> A_WL<394> A_WL<393> A_WL<392> A_WL<391> A_WL<390> A_WL<389> A_WL<388> A_WL<387> A_WL<386> A_WL<385> A_WL<384> A_WL<383> A_WL<382> A_WL<381> A_WL<380> A_WL<379> A_WL<378> A_WL<377> A_WL<376> A_WL<375> A_WL<374> A_WL<373> A_WL<372> A_WL<371> A_WL<370> A_WL<369> A_WL<368> A_WL<367> A_WL<366> A_WL<365> A_WL<364> A_WL<363> A_WL<362> A_WL<361> A_WL<360> A_WL<359> A_WL<358> A_WL<357> A_WL<356> A_WL<355> A_WL<354> A_WL<353> A_WL<352> A_WL<351> A_WL<350> A_WL<349> A_WL<348> A_WL<347> A_WL<346> A_WL<345> A_WL<344> A_WL<343> A_WL<342> A_WL<341> A_WL<340> A_WL<339> A_WL<338> A_WL<337> A_WL<336> A_WL<335> A_WL<334> A_WL<333> A_WL<332> A_WL<331> A_WL<330> A_WL<329> A_WL<328> A_WL<327> A_WL<326> A_WL<325> A_WL<324> A_WL<323> A_WL<322> A_WL<321> A_WL<320> A_WL<319> A_WL<318> A_WL<317> A_WL<316> A_WL<315> A_WL<314> A_WL<313> A_WL<312> A_WL<311> A_WL<310> A_WL<309> A_WL<308> A_WL<307> A_WL<306> A_WL<305> A_WL<304> A_WL<303> A_WL<302> A_WL<301> A_WL<300> A_WL<299> A_WL<298> A_WL<297> A_WL<296> A_WL<295> A_WL<294> A_WL<293> A_WL<292> A_WL<291> A_WL<290> A_WL<289> A_WL<288> A_WL<287> A_WL<286> A_WL<285> A_WL<284> A_WL<283> A_WL<282> A_WL<281> A_WL<280> A_WL<279> A_WL<278> A_WL<277> A_WL<276> A_WL<275> A_WL<274> A_WL<273> A_WL<272> A_WL<271> A_WL<270> A_WL<269> A_WL<268> A_WL<267> A_WL<266> A_WL<265> A_WL<264> A_WL<263> A_WL<262> A_WL<261> A_WL<260> A_WL<259> A_WL<258> A_WL<257> A_WL<256> A_WL<255> A_WL<254> A_WL<253> A_WL<252> A_WL<251> A_WL<250> A_WL<249> A_WL<248> A_WL<247> A_WL<246> A_WL<245> A_WL<244> A_WL<243> A_WL<242> A_WL<241> A_WL<240> A_WL<239> A_WL<238> A_WL<237> A_WL<236> A_WL<235> A_WL<234> A_WL<233> A_WL<232> A_WL<231> A_WL<230> A_WL<229> A_WL<228> A_WL<227> A_WL<226> A_WL<225> A_WL<224> A_WL<223> A_WL<222> A_WL<221> A_WL<220> A_WL<219> A_WL<218> A_WL<217> A_WL<216> A_WL<215> A_WL<214> A_WL<213> A_WL<212> A_WL<211> A_WL<210> A_WL<209> A_WL<208> A_WL<207> A_WL<206> A_WL<205> A_WL<204> A_WL<203> A_WL<202> A_WL<201> A_WL<200> A_WL<199> A_WL<198> A_WL<197> A_WL<196> A_WL<195> A_WL<194> A_WL<193> A_WL<192> A_WL<191> A_WL<190> A_WL<189> A_WL<188> A_WL<187> A_WL<186> A_WL<185> A_WL<184> A_WL<183> A_WL<182> A_WL<181> A_WL<180> A_WL<179> A_WL<178> A_WL<177> A_WL<176> A_WL<175> A_WL<174> A_WL<173> A_WL<172> A_WL<171> A_WL<170> A_WL<169> A_WL<168> A_WL<167> A_WL<166> A_WL<165> A_WL<164> A_WL<163> A_WL<162> A_WL<161> A_WL<160> A_WL<159> A_WL<158> A_WL<157> A_WL<156> A_WL<155> A_WL<154> A_WL<153> A_WL<152> A_WL<151> A_WL<150> A_WL<149> A_WL<148> A_WL<147> A_WL<146> A_WL<145> A_WL<144> A_WL<143> A_WL<142> A_WL<141> A_WL<140> A_WL<139> A_WL<138> A_WL<137> A_WL<136> A_WL<135> A_WL<134> A_WL<133> A_WL<132> A_WL<131> A_WL<130> A_WL<129> A_WL<128> A_WL<127> A_WL<126> A_WL<125> A_WL<124> A_WL<123> A_WL<122> A_WL<121> A_WL<120> A_WL<119> A_WL<118> A_WL<117> A_WL<116> A_WL<115> A_WL<114> A_WL<113> A_WL<112> A_WL<111> A_WL<110> A_WL<109> A_WL<108> A_WL<107> A_WL<106> A_WL<105> A_WL<104> A_WL<103> A_WL<102> A_WL<101> A_WL<100> A_WL<99> A_WL<98> A_WL<97> A_WL<96> A_WL<95> A_WL<94> A_WL<93> A_WL<92> A_WL<91> A_WL<90> A_WL<89> A_WL<88> A_WL<87> A_WL<86> A_WL<85> A_WL<84> A_WL<83> A_WL<82> A_WL<81> A_WL<80> A_WL<79> A_WL<78> A_WL<77> A_WL<76> A_WL<75> A_WL<74> A_WL<73> A_WL<72> A_WL<71> A_WL<70> A_WL<69> A_WL<68> A_WL<67> A_WL<66> A_WL<65> A_WL<64> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS
XCORNER<3> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_CORNER
XCORNER<2> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_CORNER
XCORNER<1> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_CORNER
XCORNER<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_CORNER
XRAMEDGE_L<31> A_WL<511> A_WL<510> A_WL<509> A_WL<508> A_WL<507> A_WL<506> A_WL<505> A_WL<504> A_WL<503> A_WL<502> A_WL<501> A_WL<500> A_WL<499> A_WL<498> A_WL<497> A_WL<496> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<30> A_WL<495> A_WL<494> A_WL<493> A_WL<492> A_WL<491> A_WL<490> A_WL<489> A_WL<488> A_WL<487> A_WL<486> A_WL<485> A_WL<484> A_WL<483> A_WL<482> A_WL<481> A_WL<480> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<29> A_WL<479> A_WL<478> A_WL<477> A_WL<476> A_WL<475> A_WL<474> A_WL<473> A_WL<472> A_WL<471> A_WL<470> A_WL<469> A_WL<468> A_WL<467> A_WL<466> A_WL<465> A_WL<464> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<28> A_WL<463> A_WL<462> A_WL<461> A_WL<460> A_WL<459> A_WL<458> A_WL<457> A_WL<456> A_WL<455> A_WL<454> A_WL<453> A_WL<452> A_WL<451> A_WL<450> A_WL<449> A_WL<448> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<27> A_WL<447> A_WL<446> A_WL<445> A_WL<444> A_WL<443> A_WL<442> A_WL<441> A_WL<440> A_WL<439> A_WL<438> A_WL<437> A_WL<436> A_WL<435> A_WL<434> A_WL<433> A_WL<432> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<26> A_WL<431> A_WL<430> A_WL<429> A_WL<428> A_WL<427> A_WL<426> A_WL<425> A_WL<424> A_WL<423> A_WL<422> A_WL<421> A_WL<420> A_WL<419> A_WL<418> A_WL<417> A_WL<416> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<25> A_WL<415> A_WL<414> A_WL<413> A_WL<412> A_WL<411> A_WL<410> A_WL<409> A_WL<408> A_WL<407> A_WL<406> A_WL<405> A_WL<404> A_WL<403> A_WL<402> A_WL<401> A_WL<400> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<24> A_WL<399> A_WL<398> A_WL<397> A_WL<396> A_WL<395> A_WL<394> A_WL<393> A_WL<392> A_WL<391> A_WL<390> A_WL<389> A_WL<388> A_WL<387> A_WL<386> A_WL<385> A_WL<384> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<23> A_WL<383> A_WL<382> A_WL<381> A_WL<380> A_WL<379> A_WL<378> A_WL<377> A_WL<376> A_WL<375> A_WL<374> A_WL<373> A_WL<372> A_WL<371> A_WL<370> A_WL<369> A_WL<368> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<22> A_WL<367> A_WL<366> A_WL<365> A_WL<364> A_WL<363> A_WL<362> A_WL<361> A_WL<360> A_WL<359> A_WL<358> A_WL<357> A_WL<356> A_WL<355> A_WL<354> A_WL<353> A_WL<352> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<21> A_WL<351> A_WL<350> A_WL<349> A_WL<348> A_WL<347> A_WL<346> A_WL<345> A_WL<344> A_WL<343> A_WL<342> A_WL<341> A_WL<340> A_WL<339> A_WL<338> A_WL<337> A_WL<336> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<20> A_WL<335> A_WL<334> A_WL<333> A_WL<332> A_WL<331> A_WL<330> A_WL<329> A_WL<328> A_WL<327> A_WL<326> A_WL<325> A_WL<324> A_WL<323> A_WL<322> A_WL<321> A_WL<320> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<19> A_WL<319> A_WL<318> A_WL<317> A_WL<316> A_WL<315> A_WL<314> A_WL<313> A_WL<312> A_WL<311> A_WL<310> A_WL<309> A_WL<308> A_WL<307> A_WL<306> A_WL<305> A_WL<304> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<18> A_WL<303> A_WL<302> A_WL<301> A_WL<300> A_WL<299> A_WL<298> A_WL<297> A_WL<296> A_WL<295> A_WL<294> A_WL<293> A_WL<292> A_WL<291> A_WL<290> A_WL<289> A_WL<288> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<17> A_WL<287> A_WL<286> A_WL<285> A_WL<284> A_WL<283> A_WL<282> A_WL<281> A_WL<280> A_WL<279> A_WL<278> A_WL<277> A_WL<276> A_WL<275> A_WL<274> A_WL<273> A_WL<272> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<16> A_WL<271> A_WL<270> A_WL<269> A_WL<268> A_WL<267> A_WL<266> A_WL<265> A_WL<264> A_WL<263> A_WL<262> A_WL<261> A_WL<260> A_WL<259> A_WL<258> A_WL<257> A_WL<256> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<15> A_WL<255> A_WL<254> A_WL<253> A_WL<252> A_WL<251> A_WL<250> A_WL<249> A_WL<248> A_WL<247> A_WL<246> A_WL<245> A_WL<244> A_WL<243> A_WL<242> A_WL<241> A_WL<240> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<14> A_WL<239> A_WL<238> A_WL<237> A_WL<236> A_WL<235> A_WL<234> A_WL<233> A_WL<232> A_WL<231> A_WL<230> A_WL<229> A_WL<228> A_WL<227> A_WL<226> A_WL<225> A_WL<224> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<13> A_WL<223> A_WL<222> A_WL<221> A_WL<220> A_WL<219> A_WL<218> A_WL<217> A_WL<216> A_WL<215> A_WL<214> A_WL<213> A_WL<212> A_WL<211> A_WL<210> A_WL<209> A_WL<208> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<12> A_WL<207> A_WL<206> A_WL<205> A_WL<204> A_WL<203> A_WL<202> A_WL<201> A_WL<200> A_WL<199> A_WL<198> A_WL<197> A_WL<196> A_WL<195> A_WL<194> A_WL<193> A_WL<192> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<11> A_WL<191> A_WL<190> A_WL<189> A_WL<188> A_WL<187> A_WL<186> A_WL<185> A_WL<184> A_WL<183> A_WL<182> A_WL<181> A_WL<180> A_WL<179> A_WL<178> A_WL<177> A_WL<176> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<10> A_WL<175> A_WL<174> A_WL<173> A_WL<172> A_WL<171> A_WL<170> A_WL<169> A_WL<168> A_WL<167> A_WL<166> A_WL<165> A_WL<164> A_WL<163> A_WL<162> A_WL<161> A_WL<160> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<9> A_WL<159> A_WL<158> A_WL<157> A_WL<156> A_WL<155> A_WL<154> A_WL<153> A_WL<152> A_WL<151> A_WL<150> A_WL<149> A_WL<148> A_WL<147> A_WL<146> A_WL<145> A_WL<144> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<8> A_WL<143> A_WL<142> A_WL<141> A_WL<140> A_WL<139> A_WL<138> A_WL<137> A_WL<136> A_WL<135> A_WL<134> A_WL<133> A_WL<132> A_WL<131> A_WL<130> A_WL<129> A_WL<128> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<7> A_WL<127> A_WL<126> A_WL<125> A_WL<124> A_WL<123> A_WL<122> A_WL<121> A_WL<120> A_WL<119> A_WL<118> A_WL<117> A_WL<116> A_WL<115> A_WL<114> A_WL<113> A_WL<112> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<6> A_WL<111> A_WL<110> A_WL<109> A_WL<108> A_WL<107> A_WL<106> A_WL<105> A_WL<104> A_WL<103> A_WL<102> A_WL<101> A_WL<100> A_WL<99> A_WL<98> A_WL<97> A_WL<96> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<5> A_WL<95> A_WL<94> A_WL<93> A_WL<92> A_WL<91> A_WL<90> A_WL<89> A_WL<88> A_WL<87> A_WL<86> A_WL<85> A_WL<84> A_WL<83> A_WL<82> A_WL<81> A_WL<80> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<4> A_WL<79> A_WL<78> A_WL<77> A_WL<76> A_WL<75> A_WL<74> A_WL<73> A_WL<72> A_WL<71> A_WL<70> A_WL<69> A_WL<68> A_WL<67> A_WL<66> A_WL<65> A_WL<64> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<3> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<2> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<1> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_L<0> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<31> A_IWL<32767> A_IWL<32766> A_IWL<32765> A_IWL<32764> A_IWL<32763> A_IWL<32762> A_IWL<32761> A_IWL<32760> A_IWL<32759> A_IWL<32758> A_IWL<32757> A_IWL<32756> A_IWL<32755> A_IWL<32754> A_IWL<32753> A_IWL<32752> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<30> A_IWL<32751> A_IWL<32750> A_IWL<32749> A_IWL<32748> A_IWL<32747> A_IWL<32746> A_IWL<32745> A_IWL<32744> A_IWL<32743> A_IWL<32742> A_IWL<32741> A_IWL<32740> A_IWL<32739> A_IWL<32738> A_IWL<32737> A_IWL<32736> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<29> A_IWL<32735> A_IWL<32734> A_IWL<32733> A_IWL<32732> A_IWL<32731> A_IWL<32730> A_IWL<32729> A_IWL<32728> A_IWL<32727> A_IWL<32726> A_IWL<32725> A_IWL<32724> A_IWL<32723> A_IWL<32722> A_IWL<32721> A_IWL<32720> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<28> A_IWL<32719> A_IWL<32718> A_IWL<32717> A_IWL<32716> A_IWL<32715> A_IWL<32714> A_IWL<32713> A_IWL<32712> A_IWL<32711> A_IWL<32710> A_IWL<32709> A_IWL<32708> A_IWL<32707> A_IWL<32706> A_IWL<32705> A_IWL<32704> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<27> A_IWL<32703> A_IWL<32702> A_IWL<32701> A_IWL<32700> A_IWL<32699> A_IWL<32698> A_IWL<32697> A_IWL<32696> A_IWL<32695> A_IWL<32694> A_IWL<32693> A_IWL<32692> A_IWL<32691> A_IWL<32690> A_IWL<32689> A_IWL<32688> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<26> A_IWL<32687> A_IWL<32686> A_IWL<32685> A_IWL<32684> A_IWL<32683> A_IWL<32682> A_IWL<32681> A_IWL<32680> A_IWL<32679> A_IWL<32678> A_IWL<32677> A_IWL<32676> A_IWL<32675> A_IWL<32674> A_IWL<32673> A_IWL<32672> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<25> A_IWL<32671> A_IWL<32670> A_IWL<32669> A_IWL<32668> A_IWL<32667> A_IWL<32666> A_IWL<32665> A_IWL<32664> A_IWL<32663> A_IWL<32662> A_IWL<32661> A_IWL<32660> A_IWL<32659> A_IWL<32658> A_IWL<32657> A_IWL<32656> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<24> A_IWL<32655> A_IWL<32654> A_IWL<32653> A_IWL<32652> A_IWL<32651> A_IWL<32650> A_IWL<32649> A_IWL<32648> A_IWL<32647> A_IWL<32646> A_IWL<32645> A_IWL<32644> A_IWL<32643> A_IWL<32642> A_IWL<32641> A_IWL<32640> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<23> A_IWL<32639> A_IWL<32638> A_IWL<32637> A_IWL<32636> A_IWL<32635> A_IWL<32634> A_IWL<32633> A_IWL<32632> A_IWL<32631> A_IWL<32630> A_IWL<32629> A_IWL<32628> A_IWL<32627> A_IWL<32626> A_IWL<32625> A_IWL<32624> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<22> A_IWL<32623> A_IWL<32622> A_IWL<32621> A_IWL<32620> A_IWL<32619> A_IWL<32618> A_IWL<32617> A_IWL<32616> A_IWL<32615> A_IWL<32614> A_IWL<32613> A_IWL<32612> A_IWL<32611> A_IWL<32610> A_IWL<32609> A_IWL<32608> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<21> A_IWL<32607> A_IWL<32606> A_IWL<32605> A_IWL<32604> A_IWL<32603> A_IWL<32602> A_IWL<32601> A_IWL<32600> A_IWL<32599> A_IWL<32598> A_IWL<32597> A_IWL<32596> A_IWL<32595> A_IWL<32594> A_IWL<32593> A_IWL<32592> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<20> A_IWL<32591> A_IWL<32590> A_IWL<32589> A_IWL<32588> A_IWL<32587> A_IWL<32586> A_IWL<32585> A_IWL<32584> A_IWL<32583> A_IWL<32582> A_IWL<32581> A_IWL<32580> A_IWL<32579> A_IWL<32578> A_IWL<32577> A_IWL<32576> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<19> A_IWL<32575> A_IWL<32574> A_IWL<32573> A_IWL<32572> A_IWL<32571> A_IWL<32570> A_IWL<32569> A_IWL<32568> A_IWL<32567> A_IWL<32566> A_IWL<32565> A_IWL<32564> A_IWL<32563> A_IWL<32562> A_IWL<32561> A_IWL<32560> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<18> A_IWL<32559> A_IWL<32558> A_IWL<32557> A_IWL<32556> A_IWL<32555> A_IWL<32554> A_IWL<32553> A_IWL<32552> A_IWL<32551> A_IWL<32550> A_IWL<32549> A_IWL<32548> A_IWL<32547> A_IWL<32546> A_IWL<32545> A_IWL<32544> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<17> A_IWL<32543> A_IWL<32542> A_IWL<32541> A_IWL<32540> A_IWL<32539> A_IWL<32538> A_IWL<32537> A_IWL<32536> A_IWL<32535> A_IWL<32534> A_IWL<32533> A_IWL<32532> A_IWL<32531> A_IWL<32530> A_IWL<32529> A_IWL<32528> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<16> A_IWL<32527> A_IWL<32526> A_IWL<32525> A_IWL<32524> A_IWL<32523> A_IWL<32522> A_IWL<32521> A_IWL<32520> A_IWL<32519> A_IWL<32518> A_IWL<32517> A_IWL<32516> A_IWL<32515> A_IWL<32514> A_IWL<32513> A_IWL<32512> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<15> A_IWL<32511> A_IWL<32510> A_IWL<32509> A_IWL<32508> A_IWL<32507> A_IWL<32506> A_IWL<32505> A_IWL<32504> A_IWL<32503> A_IWL<32502> A_IWL<32501> A_IWL<32500> A_IWL<32499> A_IWL<32498> A_IWL<32497> A_IWL<32496> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<14> A_IWL<32495> A_IWL<32494> A_IWL<32493> A_IWL<32492> A_IWL<32491> A_IWL<32490> A_IWL<32489> A_IWL<32488> A_IWL<32487> A_IWL<32486> A_IWL<32485> A_IWL<32484> A_IWL<32483> A_IWL<32482> A_IWL<32481> A_IWL<32480> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<13> A_IWL<32479> A_IWL<32478> A_IWL<32477> A_IWL<32476> A_IWL<32475> A_IWL<32474> A_IWL<32473> A_IWL<32472> A_IWL<32471> A_IWL<32470> A_IWL<32469> A_IWL<32468> A_IWL<32467> A_IWL<32466> A_IWL<32465> A_IWL<32464> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<12> A_IWL<32463> A_IWL<32462> A_IWL<32461> A_IWL<32460> A_IWL<32459> A_IWL<32458> A_IWL<32457> A_IWL<32456> A_IWL<32455> A_IWL<32454> A_IWL<32453> A_IWL<32452> A_IWL<32451> A_IWL<32450> A_IWL<32449> A_IWL<32448> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<11> A_IWL<32447> A_IWL<32446> A_IWL<32445> A_IWL<32444> A_IWL<32443> A_IWL<32442> A_IWL<32441> A_IWL<32440> A_IWL<32439> A_IWL<32438> A_IWL<32437> A_IWL<32436> A_IWL<32435> A_IWL<32434> A_IWL<32433> A_IWL<32432> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<10> A_IWL<32431> A_IWL<32430> A_IWL<32429> A_IWL<32428> A_IWL<32427> A_IWL<32426> A_IWL<32425> A_IWL<32424> A_IWL<32423> A_IWL<32422> A_IWL<32421> A_IWL<32420> A_IWL<32419> A_IWL<32418> A_IWL<32417> A_IWL<32416> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<9> A_IWL<32415> A_IWL<32414> A_IWL<32413> A_IWL<32412> A_IWL<32411> A_IWL<32410> A_IWL<32409> A_IWL<32408> A_IWL<32407> A_IWL<32406> A_IWL<32405> A_IWL<32404> A_IWL<32403> A_IWL<32402> A_IWL<32401> A_IWL<32400> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<8> A_IWL<32399> A_IWL<32398> A_IWL<32397> A_IWL<32396> A_IWL<32395> A_IWL<32394> A_IWL<32393> A_IWL<32392> A_IWL<32391> A_IWL<32390> A_IWL<32389> A_IWL<32388> A_IWL<32387> A_IWL<32386> A_IWL<32385> A_IWL<32384> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<7> A_IWL<32383> A_IWL<32382> A_IWL<32381> A_IWL<32380> A_IWL<32379> A_IWL<32378> A_IWL<32377> A_IWL<32376> A_IWL<32375> A_IWL<32374> A_IWL<32373> A_IWL<32372> A_IWL<32371> A_IWL<32370> A_IWL<32369> A_IWL<32368> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<6> A_IWL<32367> A_IWL<32366> A_IWL<32365> A_IWL<32364> A_IWL<32363> A_IWL<32362> A_IWL<32361> A_IWL<32360> A_IWL<32359> A_IWL<32358> A_IWL<32357> A_IWL<32356> A_IWL<32355> A_IWL<32354> A_IWL<32353> A_IWL<32352> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<5> A_IWL<32351> A_IWL<32350> A_IWL<32349> A_IWL<32348> A_IWL<32347> A_IWL<32346> A_IWL<32345> A_IWL<32344> A_IWL<32343> A_IWL<32342> A_IWL<32341> A_IWL<32340> A_IWL<32339> A_IWL<32338> A_IWL<32337> A_IWL<32336> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<4> A_IWL<32335> A_IWL<32334> A_IWL<32333> A_IWL<32332> A_IWL<32331> A_IWL<32330> A_IWL<32329> A_IWL<32328> A_IWL<32327> A_IWL<32326> A_IWL<32325> A_IWL<32324> A_IWL<32323> A_IWL<32322> A_IWL<32321> A_IWL<32320> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<3> A_IWL<32319> A_IWL<32318> A_IWL<32317> A_IWL<32316> A_IWL<32315> A_IWL<32314> A_IWL<32313> A_IWL<32312> A_IWL<32311> A_IWL<32310> A_IWL<32309> A_IWL<32308> A_IWL<32307> A_IWL<32306> A_IWL<32305> A_IWL<32304> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<2> A_IWL<32303> A_IWL<32302> A_IWL<32301> A_IWL<32300> A_IWL<32299> A_IWL<32298> A_IWL<32297> A_IWL<32296> A_IWL<32295> A_IWL<32294> A_IWL<32293> A_IWL<32292> A_IWL<32291> A_IWL<32290> A_IWL<32289> A_IWL<32288> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<1> A_IWL<32287> A_IWL<32286> A_IWL<32285> A_IWL<32284> A_IWL<32283> A_IWL<32282> A_IWL<32281> A_IWL<32280> A_IWL<32279> A_IWL<32278> A_IWL<32277> A_IWL<32276> A_IWL<32275> A_IWL<32274> A_IWL<32273> A_IWL<32272> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XRAMEDGE_R<0> A_IWL<32271> A_IWL<32270> A_IWL<32269> A_IWL<32268> A_IWL<32267> A_IWL<32266> A_IWL<32265> A_IWL<32264> A_IWL<32263> A_IWL<32262> A_IWL<32261> A_IWL<32260> A_IWL<32259> A_IWL<32258> A_IWL<32257> A_IWL<32256> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_BITKIT_16x2_EDGE_LR
XCOL<63> A_BLC<127> A_BLC<126> A_BLC_TOP<127> A_BLC_TOP<126> A_BLT<127> A_BLT<126> A_BLT_TOP<127> A_BLT_TOP<126> A_IWL<32255> A_IWL<32254> A_IWL<32253> A_IWL<32252> A_IWL<32251> A_IWL<32250> A_IWL<32249> A_IWL<32248> A_IWL<32247> A_IWL<32246> A_IWL<32245> A_IWL<32244> A_IWL<32243> A_IWL<32242> A_IWL<32241> A_IWL<32240> A_IWL<32239> A_IWL<32238> A_IWL<32237> A_IWL<32236> A_IWL<32235> A_IWL<32234> A_IWL<32233> A_IWL<32232> A_IWL<32231> A_IWL<32230> A_IWL<32229> A_IWL<32228> A_IWL<32227> A_IWL<32226> A_IWL<32225> A_IWL<32224> A_IWL<32223> A_IWL<32222> A_IWL<32221> A_IWL<32220> A_IWL<32219> A_IWL<32218> A_IWL<32217> A_IWL<32216> A_IWL<32215> A_IWL<32214> A_IWL<32213> A_IWL<32212> A_IWL<32211> A_IWL<32210> A_IWL<32209> A_IWL<32208> A_IWL<32207> A_IWL<32206> A_IWL<32205> A_IWL<32204> A_IWL<32203> A_IWL<32202> A_IWL<32201> A_IWL<32200> A_IWL<32199> A_IWL<32198> A_IWL<32197> A_IWL<32196> A_IWL<32195> A_IWL<32194> A_IWL<32193> A_IWL<32192> A_IWL<32191> A_IWL<32190> A_IWL<32189> A_IWL<32188> A_IWL<32187> A_IWL<32186> A_IWL<32185> A_IWL<32184> A_IWL<32183> A_IWL<32182> A_IWL<32181> A_IWL<32180> A_IWL<32179> A_IWL<32178> A_IWL<32177> A_IWL<32176> A_IWL<32175> A_IWL<32174> A_IWL<32173> A_IWL<32172> A_IWL<32171> A_IWL<32170> A_IWL<32169> A_IWL<32168> A_IWL<32167> A_IWL<32166> A_IWL<32165> A_IWL<32164> A_IWL<32163> A_IWL<32162> A_IWL<32161> A_IWL<32160> A_IWL<32159> A_IWL<32158> A_IWL<32157> A_IWL<32156> A_IWL<32155> A_IWL<32154> A_IWL<32153> A_IWL<32152> A_IWL<32151> A_IWL<32150> A_IWL<32149> A_IWL<32148> A_IWL<32147> A_IWL<32146> A_IWL<32145> A_IWL<32144> A_IWL<32143> A_IWL<32142> A_IWL<32141> A_IWL<32140> A_IWL<32139> A_IWL<32138> A_IWL<32137> A_IWL<32136> A_IWL<32135> A_IWL<32134> A_IWL<32133> A_IWL<32132> A_IWL<32131> A_IWL<32130> A_IWL<32129> A_IWL<32128> A_IWL<32127> A_IWL<32126> A_IWL<32125> A_IWL<32124> A_IWL<32123> A_IWL<32122> A_IWL<32121> A_IWL<32120> A_IWL<32119> A_IWL<32118> A_IWL<32117> A_IWL<32116> A_IWL<32115> A_IWL<32114> A_IWL<32113> A_IWL<32112> A_IWL<32111> A_IWL<32110> A_IWL<32109> A_IWL<32108> A_IWL<32107> A_IWL<32106> A_IWL<32105> A_IWL<32104> A_IWL<32103> A_IWL<32102> A_IWL<32101> A_IWL<32100> A_IWL<32099> A_IWL<32098> A_IWL<32097> A_IWL<32096> A_IWL<32095> A_IWL<32094> A_IWL<32093> A_IWL<32092> A_IWL<32091> A_IWL<32090> A_IWL<32089> A_IWL<32088> A_IWL<32087> A_IWL<32086> A_IWL<32085> A_IWL<32084> A_IWL<32083> A_IWL<32082> A_IWL<32081> A_IWL<32080> A_IWL<32079> A_IWL<32078> A_IWL<32077> A_IWL<32076> A_IWL<32075> A_IWL<32074> A_IWL<32073> A_IWL<32072> A_IWL<32071> A_IWL<32070> A_IWL<32069> A_IWL<32068> A_IWL<32067> A_IWL<32066> A_IWL<32065> A_IWL<32064> A_IWL<32063> A_IWL<32062> A_IWL<32061> A_IWL<32060> A_IWL<32059> A_IWL<32058> A_IWL<32057> A_IWL<32056> A_IWL<32055> A_IWL<32054> A_IWL<32053> A_IWL<32052> A_IWL<32051> A_IWL<32050> A_IWL<32049> A_IWL<32048> A_IWL<32047> A_IWL<32046> A_IWL<32045> A_IWL<32044> A_IWL<32043> A_IWL<32042> A_IWL<32041> A_IWL<32040> A_IWL<32039> A_IWL<32038> A_IWL<32037> A_IWL<32036> A_IWL<32035> A_IWL<32034> A_IWL<32033> A_IWL<32032> A_IWL<32031> A_IWL<32030> A_IWL<32029> A_IWL<32028> A_IWL<32027> A_IWL<32026> A_IWL<32025> A_IWL<32024> A_IWL<32023> A_IWL<32022> A_IWL<32021> A_IWL<32020> A_IWL<32019> A_IWL<32018> A_IWL<32017> A_IWL<32016> A_IWL<32015> A_IWL<32014> A_IWL<32013> A_IWL<32012> A_IWL<32011> A_IWL<32010> A_IWL<32009> A_IWL<32008> A_IWL<32007> A_IWL<32006> A_IWL<32005> A_IWL<32004> A_IWL<32003> A_IWL<32002> A_IWL<32001> A_IWL<32000> A_IWL<31999> A_IWL<31998> A_IWL<31997> A_IWL<31996> A_IWL<31995> A_IWL<31994> A_IWL<31993> A_IWL<31992> A_IWL<31991> A_IWL<31990> A_IWL<31989> A_IWL<31988> A_IWL<31987> A_IWL<31986> A_IWL<31985> A_IWL<31984> A_IWL<31983> A_IWL<31982> A_IWL<31981> A_IWL<31980> A_IWL<31979> A_IWL<31978> A_IWL<31977> A_IWL<31976> A_IWL<31975> A_IWL<31974> A_IWL<31973> A_IWL<31972> A_IWL<31971> A_IWL<31970> A_IWL<31969> A_IWL<31968> A_IWL<31967> A_IWL<31966> A_IWL<31965> A_IWL<31964> A_IWL<31963> A_IWL<31962> A_IWL<31961> A_IWL<31960> A_IWL<31959> A_IWL<31958> A_IWL<31957> A_IWL<31956> A_IWL<31955> A_IWL<31954> A_IWL<31953> A_IWL<31952> A_IWL<31951> A_IWL<31950> A_IWL<31949> A_IWL<31948> A_IWL<31947> A_IWL<31946> A_IWL<31945> A_IWL<31944> A_IWL<31943> A_IWL<31942> A_IWL<31941> A_IWL<31940> A_IWL<31939> A_IWL<31938> A_IWL<31937> A_IWL<31936> A_IWL<31935> A_IWL<31934> A_IWL<31933> A_IWL<31932> A_IWL<31931> A_IWL<31930> A_IWL<31929> A_IWL<31928> A_IWL<31927> A_IWL<31926> A_IWL<31925> A_IWL<31924> A_IWL<31923> A_IWL<31922> A_IWL<31921> A_IWL<31920> A_IWL<31919> A_IWL<31918> A_IWL<31917> A_IWL<31916> A_IWL<31915> A_IWL<31914> A_IWL<31913> A_IWL<31912> A_IWL<31911> A_IWL<31910> A_IWL<31909> A_IWL<31908> A_IWL<31907> A_IWL<31906> A_IWL<31905> A_IWL<31904> A_IWL<31903> A_IWL<31902> A_IWL<31901> A_IWL<31900> A_IWL<31899> A_IWL<31898> A_IWL<31897> A_IWL<31896> A_IWL<31895> A_IWL<31894> A_IWL<31893> A_IWL<31892> A_IWL<31891> A_IWL<31890> A_IWL<31889> A_IWL<31888> A_IWL<31887> A_IWL<31886> A_IWL<31885> A_IWL<31884> A_IWL<31883> A_IWL<31882> A_IWL<31881> A_IWL<31880> A_IWL<31879> A_IWL<31878> A_IWL<31877> A_IWL<31876> A_IWL<31875> A_IWL<31874> A_IWL<31873> A_IWL<31872> A_IWL<31871> A_IWL<31870> A_IWL<31869> A_IWL<31868> A_IWL<31867> A_IWL<31866> A_IWL<31865> A_IWL<31864> A_IWL<31863> A_IWL<31862> A_IWL<31861> A_IWL<31860> A_IWL<31859> A_IWL<31858> A_IWL<31857> A_IWL<31856> A_IWL<31855> A_IWL<31854> A_IWL<31853> A_IWL<31852> A_IWL<31851> A_IWL<31850> A_IWL<31849> A_IWL<31848> A_IWL<31847> A_IWL<31846> A_IWL<31845> A_IWL<31844> A_IWL<31843> A_IWL<31842> A_IWL<31841> A_IWL<31840> A_IWL<31839> A_IWL<31838> A_IWL<31837> A_IWL<31836> A_IWL<31835> A_IWL<31834> A_IWL<31833> A_IWL<31832> A_IWL<31831> A_IWL<31830> A_IWL<31829> A_IWL<31828> A_IWL<31827> A_IWL<31826> A_IWL<31825> A_IWL<31824> A_IWL<31823> A_IWL<31822> A_IWL<31821> A_IWL<31820> A_IWL<31819> A_IWL<31818> A_IWL<31817> A_IWL<31816> A_IWL<31815> A_IWL<31814> A_IWL<31813> A_IWL<31812> A_IWL<31811> A_IWL<31810> A_IWL<31809> A_IWL<31808> A_IWL<31807> A_IWL<31806> A_IWL<31805> A_IWL<31804> A_IWL<31803> A_IWL<31802> A_IWL<31801> A_IWL<31800> A_IWL<31799> A_IWL<31798> A_IWL<31797> A_IWL<31796> A_IWL<31795> A_IWL<31794> A_IWL<31793> A_IWL<31792> A_IWL<31791> A_IWL<31790> A_IWL<31789> A_IWL<31788> A_IWL<31787> A_IWL<31786> A_IWL<31785> A_IWL<31784> A_IWL<31783> A_IWL<31782> A_IWL<31781> A_IWL<31780> A_IWL<31779> A_IWL<31778> A_IWL<31777> A_IWL<31776> A_IWL<31775> A_IWL<31774> A_IWL<31773> A_IWL<31772> A_IWL<31771> A_IWL<31770> A_IWL<31769> A_IWL<31768> A_IWL<31767> A_IWL<31766> A_IWL<31765> A_IWL<31764> A_IWL<31763> A_IWL<31762> A_IWL<31761> A_IWL<31760> A_IWL<31759> A_IWL<31758> A_IWL<31757> A_IWL<31756> A_IWL<31755> A_IWL<31754> A_IWL<31753> A_IWL<31752> A_IWL<31751> A_IWL<31750> A_IWL<31749> A_IWL<31748> A_IWL<31747> A_IWL<31746> A_IWL<31745> A_IWL<31744> A_IWL<32767> A_IWL<32766> A_IWL<32765> A_IWL<32764> A_IWL<32763> A_IWL<32762> A_IWL<32761> A_IWL<32760> A_IWL<32759> A_IWL<32758> A_IWL<32757> A_IWL<32756> A_IWL<32755> A_IWL<32754> A_IWL<32753> A_IWL<32752> A_IWL<32751> A_IWL<32750> A_IWL<32749> A_IWL<32748> A_IWL<32747> A_IWL<32746> A_IWL<32745> A_IWL<32744> A_IWL<32743> A_IWL<32742> A_IWL<32741> A_IWL<32740> A_IWL<32739> A_IWL<32738> A_IWL<32737> A_IWL<32736> A_IWL<32735> A_IWL<32734> A_IWL<32733> A_IWL<32732> A_IWL<32731> A_IWL<32730> A_IWL<32729> A_IWL<32728> A_IWL<32727> A_IWL<32726> A_IWL<32725> A_IWL<32724> A_IWL<32723> A_IWL<32722> A_IWL<32721> A_IWL<32720> A_IWL<32719> A_IWL<32718> A_IWL<32717> A_IWL<32716> A_IWL<32715> A_IWL<32714> A_IWL<32713> A_IWL<32712> A_IWL<32711> A_IWL<32710> A_IWL<32709> A_IWL<32708> A_IWL<32707> A_IWL<32706> A_IWL<32705> A_IWL<32704> A_IWL<32703> A_IWL<32702> A_IWL<32701> A_IWL<32700> A_IWL<32699> A_IWL<32698> A_IWL<32697> A_IWL<32696> A_IWL<32695> A_IWL<32694> A_IWL<32693> A_IWL<32692> A_IWL<32691> A_IWL<32690> A_IWL<32689> A_IWL<32688> A_IWL<32687> A_IWL<32686> A_IWL<32685> A_IWL<32684> A_IWL<32683> A_IWL<32682> A_IWL<32681> A_IWL<32680> A_IWL<32679> A_IWL<32678> A_IWL<32677> A_IWL<32676> A_IWL<32675> A_IWL<32674> A_IWL<32673> A_IWL<32672> A_IWL<32671> A_IWL<32670> A_IWL<32669> A_IWL<32668> A_IWL<32667> A_IWL<32666> A_IWL<32665> A_IWL<32664> A_IWL<32663> A_IWL<32662> A_IWL<32661> A_IWL<32660> A_IWL<32659> A_IWL<32658> A_IWL<32657> A_IWL<32656> A_IWL<32655> A_IWL<32654> A_IWL<32653> A_IWL<32652> A_IWL<32651> A_IWL<32650> A_IWL<32649> A_IWL<32648> A_IWL<32647> A_IWL<32646> A_IWL<32645> A_IWL<32644> A_IWL<32643> A_IWL<32642> A_IWL<32641> A_IWL<32640> A_IWL<32639> A_IWL<32638> A_IWL<32637> A_IWL<32636> A_IWL<32635> A_IWL<32634> A_IWL<32633> A_IWL<32632> A_IWL<32631> A_IWL<32630> A_IWL<32629> A_IWL<32628> A_IWL<32627> A_IWL<32626> A_IWL<32625> A_IWL<32624> A_IWL<32623> A_IWL<32622> A_IWL<32621> A_IWL<32620> A_IWL<32619> A_IWL<32618> A_IWL<32617> A_IWL<32616> A_IWL<32615> A_IWL<32614> A_IWL<32613> A_IWL<32612> A_IWL<32611> A_IWL<32610> A_IWL<32609> A_IWL<32608> A_IWL<32607> A_IWL<32606> A_IWL<32605> A_IWL<32604> A_IWL<32603> A_IWL<32602> A_IWL<32601> A_IWL<32600> A_IWL<32599> A_IWL<32598> A_IWL<32597> A_IWL<32596> A_IWL<32595> A_IWL<32594> A_IWL<32593> A_IWL<32592> A_IWL<32591> A_IWL<32590> A_IWL<32589> A_IWL<32588> A_IWL<32587> A_IWL<32586> A_IWL<32585> A_IWL<32584> A_IWL<32583> A_IWL<32582> A_IWL<32581> A_IWL<32580> A_IWL<32579> A_IWL<32578> A_IWL<32577> A_IWL<32576> A_IWL<32575> A_IWL<32574> A_IWL<32573> A_IWL<32572> A_IWL<32571> A_IWL<32570> A_IWL<32569> A_IWL<32568> A_IWL<32567> A_IWL<32566> A_IWL<32565> A_IWL<32564> A_IWL<32563> A_IWL<32562> A_IWL<32561> A_IWL<32560> A_IWL<32559> A_IWL<32558> A_IWL<32557> A_IWL<32556> A_IWL<32555> A_IWL<32554> A_IWL<32553> A_IWL<32552> A_IWL<32551> A_IWL<32550> A_IWL<32549> A_IWL<32548> A_IWL<32547> A_IWL<32546> A_IWL<32545> A_IWL<32544> A_IWL<32543> A_IWL<32542> A_IWL<32541> A_IWL<32540> A_IWL<32539> A_IWL<32538> A_IWL<32537> A_IWL<32536> A_IWL<32535> A_IWL<32534> A_IWL<32533> A_IWL<32532> A_IWL<32531> A_IWL<32530> A_IWL<32529> A_IWL<32528> A_IWL<32527> A_IWL<32526> A_IWL<32525> A_IWL<32524> A_IWL<32523> A_IWL<32522> A_IWL<32521> A_IWL<32520> A_IWL<32519> A_IWL<32518> A_IWL<32517> A_IWL<32516> A_IWL<32515> A_IWL<32514> A_IWL<32513> A_IWL<32512> A_IWL<32511> A_IWL<32510> A_IWL<32509> A_IWL<32508> A_IWL<32507> A_IWL<32506> A_IWL<32505> A_IWL<32504> A_IWL<32503> A_IWL<32502> A_IWL<32501> A_IWL<32500> A_IWL<32499> A_IWL<32498> A_IWL<32497> A_IWL<32496> A_IWL<32495> A_IWL<32494> A_IWL<32493> A_IWL<32492> A_IWL<32491> A_IWL<32490> A_IWL<32489> A_IWL<32488> A_IWL<32487> A_IWL<32486> A_IWL<32485> A_IWL<32484> A_IWL<32483> A_IWL<32482> A_IWL<32481> A_IWL<32480> A_IWL<32479> A_IWL<32478> A_IWL<32477> A_IWL<32476> A_IWL<32475> A_IWL<32474> A_IWL<32473> A_IWL<32472> A_IWL<32471> A_IWL<32470> A_IWL<32469> A_IWL<32468> A_IWL<32467> A_IWL<32466> A_IWL<32465> A_IWL<32464> A_IWL<32463> A_IWL<32462> A_IWL<32461> A_IWL<32460> A_IWL<32459> A_IWL<32458> A_IWL<32457> A_IWL<32456> A_IWL<32455> A_IWL<32454> A_IWL<32453> A_IWL<32452> A_IWL<32451> A_IWL<32450> A_IWL<32449> A_IWL<32448> A_IWL<32447> A_IWL<32446> A_IWL<32445> A_IWL<32444> A_IWL<32443> A_IWL<32442> A_IWL<32441> A_IWL<32440> A_IWL<32439> A_IWL<32438> A_IWL<32437> A_IWL<32436> A_IWL<32435> A_IWL<32434> A_IWL<32433> A_IWL<32432> A_IWL<32431> A_IWL<32430> A_IWL<32429> A_IWL<32428> A_IWL<32427> A_IWL<32426> A_IWL<32425> A_IWL<32424> A_IWL<32423> A_IWL<32422> A_IWL<32421> A_IWL<32420> A_IWL<32419> A_IWL<32418> A_IWL<32417> A_IWL<32416> A_IWL<32415> A_IWL<32414> A_IWL<32413> A_IWL<32412> A_IWL<32411> A_IWL<32410> A_IWL<32409> A_IWL<32408> A_IWL<32407> A_IWL<32406> A_IWL<32405> A_IWL<32404> A_IWL<32403> A_IWL<32402> A_IWL<32401> A_IWL<32400> A_IWL<32399> A_IWL<32398> A_IWL<32397> A_IWL<32396> A_IWL<32395> A_IWL<32394> A_IWL<32393> A_IWL<32392> A_IWL<32391> A_IWL<32390> A_IWL<32389> A_IWL<32388> A_IWL<32387> A_IWL<32386> A_IWL<32385> A_IWL<32384> A_IWL<32383> A_IWL<32382> A_IWL<32381> A_IWL<32380> A_IWL<32379> A_IWL<32378> A_IWL<32377> A_IWL<32376> A_IWL<32375> A_IWL<32374> A_IWL<32373> A_IWL<32372> A_IWL<32371> A_IWL<32370> A_IWL<32369> A_IWL<32368> A_IWL<32367> A_IWL<32366> A_IWL<32365> A_IWL<32364> A_IWL<32363> A_IWL<32362> A_IWL<32361> A_IWL<32360> A_IWL<32359> A_IWL<32358> A_IWL<32357> A_IWL<32356> A_IWL<32355> A_IWL<32354> A_IWL<32353> A_IWL<32352> A_IWL<32351> A_IWL<32350> A_IWL<32349> A_IWL<32348> A_IWL<32347> A_IWL<32346> A_IWL<32345> A_IWL<32344> A_IWL<32343> A_IWL<32342> A_IWL<32341> A_IWL<32340> A_IWL<32339> A_IWL<32338> A_IWL<32337> A_IWL<32336> A_IWL<32335> A_IWL<32334> A_IWL<32333> A_IWL<32332> A_IWL<32331> A_IWL<32330> A_IWL<32329> A_IWL<32328> A_IWL<32327> A_IWL<32326> A_IWL<32325> A_IWL<32324> A_IWL<32323> A_IWL<32322> A_IWL<32321> A_IWL<32320> A_IWL<32319> A_IWL<32318> A_IWL<32317> A_IWL<32316> A_IWL<32315> A_IWL<32314> A_IWL<32313> A_IWL<32312> A_IWL<32311> A_IWL<32310> A_IWL<32309> A_IWL<32308> A_IWL<32307> A_IWL<32306> A_IWL<32305> A_IWL<32304> A_IWL<32303> A_IWL<32302> A_IWL<32301> A_IWL<32300> A_IWL<32299> A_IWL<32298> A_IWL<32297> A_IWL<32296> A_IWL<32295> A_IWL<32294> A_IWL<32293> A_IWL<32292> A_IWL<32291> A_IWL<32290> A_IWL<32289> A_IWL<32288> A_IWL<32287> A_IWL<32286> A_IWL<32285> A_IWL<32284> A_IWL<32283> A_IWL<32282> A_IWL<32281> A_IWL<32280> A_IWL<32279> A_IWL<32278> A_IWL<32277> A_IWL<32276> A_IWL<32275> A_IWL<32274> A_IWL<32273> A_IWL<32272> A_IWL<32271> A_IWL<32270> A_IWL<32269> A_IWL<32268> A_IWL<32267> A_IWL<32266> A_IWL<32265> A_IWL<32264> A_IWL<32263> A_IWL<32262> A_IWL<32261> A_IWL<32260> A_IWL<32259> A_IWL<32258> A_IWL<32257> A_IWL<32256> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<62> A_BLC<125> A_BLC<124> A_BLC_TOP<125> A_BLC_TOP<124> A_BLT<125> A_BLT<124> A_BLT_TOP<125> A_BLT_TOP<124> A_IWL<31743> A_IWL<31742> A_IWL<31741> A_IWL<31740> A_IWL<31739> A_IWL<31738> A_IWL<31737> A_IWL<31736> A_IWL<31735> A_IWL<31734> A_IWL<31733> A_IWL<31732> A_IWL<31731> A_IWL<31730> A_IWL<31729> A_IWL<31728> A_IWL<31727> A_IWL<31726> A_IWL<31725> A_IWL<31724> A_IWL<31723> A_IWL<31722> A_IWL<31721> A_IWL<31720> A_IWL<31719> A_IWL<31718> A_IWL<31717> A_IWL<31716> A_IWL<31715> A_IWL<31714> A_IWL<31713> A_IWL<31712> A_IWL<31711> A_IWL<31710> A_IWL<31709> A_IWL<31708> A_IWL<31707> A_IWL<31706> A_IWL<31705> A_IWL<31704> A_IWL<31703> A_IWL<31702> A_IWL<31701> A_IWL<31700> A_IWL<31699> A_IWL<31698> A_IWL<31697> A_IWL<31696> A_IWL<31695> A_IWL<31694> A_IWL<31693> A_IWL<31692> A_IWL<31691> A_IWL<31690> A_IWL<31689> A_IWL<31688> A_IWL<31687> A_IWL<31686> A_IWL<31685> A_IWL<31684> A_IWL<31683> A_IWL<31682> A_IWL<31681> A_IWL<31680> A_IWL<31679> A_IWL<31678> A_IWL<31677> A_IWL<31676> A_IWL<31675> A_IWL<31674> A_IWL<31673> A_IWL<31672> A_IWL<31671> A_IWL<31670> A_IWL<31669> A_IWL<31668> A_IWL<31667> A_IWL<31666> A_IWL<31665> A_IWL<31664> A_IWL<31663> A_IWL<31662> A_IWL<31661> A_IWL<31660> A_IWL<31659> A_IWL<31658> A_IWL<31657> A_IWL<31656> A_IWL<31655> A_IWL<31654> A_IWL<31653> A_IWL<31652> A_IWL<31651> A_IWL<31650> A_IWL<31649> A_IWL<31648> A_IWL<31647> A_IWL<31646> A_IWL<31645> A_IWL<31644> A_IWL<31643> A_IWL<31642> A_IWL<31641> A_IWL<31640> A_IWL<31639> A_IWL<31638> A_IWL<31637> A_IWL<31636> A_IWL<31635> A_IWL<31634> A_IWL<31633> A_IWL<31632> A_IWL<31631> A_IWL<31630> A_IWL<31629> A_IWL<31628> A_IWL<31627> A_IWL<31626> A_IWL<31625> A_IWL<31624> A_IWL<31623> A_IWL<31622> A_IWL<31621> A_IWL<31620> A_IWL<31619> A_IWL<31618> A_IWL<31617> A_IWL<31616> A_IWL<31615> A_IWL<31614> A_IWL<31613> A_IWL<31612> A_IWL<31611> A_IWL<31610> A_IWL<31609> A_IWL<31608> A_IWL<31607> A_IWL<31606> A_IWL<31605> A_IWL<31604> A_IWL<31603> A_IWL<31602> A_IWL<31601> A_IWL<31600> A_IWL<31599> A_IWL<31598> A_IWL<31597> A_IWL<31596> A_IWL<31595> A_IWL<31594> A_IWL<31593> A_IWL<31592> A_IWL<31591> A_IWL<31590> A_IWL<31589> A_IWL<31588> A_IWL<31587> A_IWL<31586> A_IWL<31585> A_IWL<31584> A_IWL<31583> A_IWL<31582> A_IWL<31581> A_IWL<31580> A_IWL<31579> A_IWL<31578> A_IWL<31577> A_IWL<31576> A_IWL<31575> A_IWL<31574> A_IWL<31573> A_IWL<31572> A_IWL<31571> A_IWL<31570> A_IWL<31569> A_IWL<31568> A_IWL<31567> A_IWL<31566> A_IWL<31565> A_IWL<31564> A_IWL<31563> A_IWL<31562> A_IWL<31561> A_IWL<31560> A_IWL<31559> A_IWL<31558> A_IWL<31557> A_IWL<31556> A_IWL<31555> A_IWL<31554> A_IWL<31553> A_IWL<31552> A_IWL<31551> A_IWL<31550> A_IWL<31549> A_IWL<31548> A_IWL<31547> A_IWL<31546> A_IWL<31545> A_IWL<31544> A_IWL<31543> A_IWL<31542> A_IWL<31541> A_IWL<31540> A_IWL<31539> A_IWL<31538> A_IWL<31537> A_IWL<31536> A_IWL<31535> A_IWL<31534> A_IWL<31533> A_IWL<31532> A_IWL<31531> A_IWL<31530> A_IWL<31529> A_IWL<31528> A_IWL<31527> A_IWL<31526> A_IWL<31525> A_IWL<31524> A_IWL<31523> A_IWL<31522> A_IWL<31521> A_IWL<31520> A_IWL<31519> A_IWL<31518> A_IWL<31517> A_IWL<31516> A_IWL<31515> A_IWL<31514> A_IWL<31513> A_IWL<31512> A_IWL<31511> A_IWL<31510> A_IWL<31509> A_IWL<31508> A_IWL<31507> A_IWL<31506> A_IWL<31505> A_IWL<31504> A_IWL<31503> A_IWL<31502> A_IWL<31501> A_IWL<31500> A_IWL<31499> A_IWL<31498> A_IWL<31497> A_IWL<31496> A_IWL<31495> A_IWL<31494> A_IWL<31493> A_IWL<31492> A_IWL<31491> A_IWL<31490> A_IWL<31489> A_IWL<31488> A_IWL<31487> A_IWL<31486> A_IWL<31485> A_IWL<31484> A_IWL<31483> A_IWL<31482> A_IWL<31481> A_IWL<31480> A_IWL<31479> A_IWL<31478> A_IWL<31477> A_IWL<31476> A_IWL<31475> A_IWL<31474> A_IWL<31473> A_IWL<31472> A_IWL<31471> A_IWL<31470> A_IWL<31469> A_IWL<31468> A_IWL<31467> A_IWL<31466> A_IWL<31465> A_IWL<31464> A_IWL<31463> A_IWL<31462> A_IWL<31461> A_IWL<31460> A_IWL<31459> A_IWL<31458> A_IWL<31457> A_IWL<31456> A_IWL<31455> A_IWL<31454> A_IWL<31453> A_IWL<31452> A_IWL<31451> A_IWL<31450> A_IWL<31449> A_IWL<31448> A_IWL<31447> A_IWL<31446> A_IWL<31445> A_IWL<31444> A_IWL<31443> A_IWL<31442> A_IWL<31441> A_IWL<31440> A_IWL<31439> A_IWL<31438> A_IWL<31437> A_IWL<31436> A_IWL<31435> A_IWL<31434> A_IWL<31433> A_IWL<31432> A_IWL<31431> A_IWL<31430> A_IWL<31429> A_IWL<31428> A_IWL<31427> A_IWL<31426> A_IWL<31425> A_IWL<31424> A_IWL<31423> A_IWL<31422> A_IWL<31421> A_IWL<31420> A_IWL<31419> A_IWL<31418> A_IWL<31417> A_IWL<31416> A_IWL<31415> A_IWL<31414> A_IWL<31413> A_IWL<31412> A_IWL<31411> A_IWL<31410> A_IWL<31409> A_IWL<31408> A_IWL<31407> A_IWL<31406> A_IWL<31405> A_IWL<31404> A_IWL<31403> A_IWL<31402> A_IWL<31401> A_IWL<31400> A_IWL<31399> A_IWL<31398> A_IWL<31397> A_IWL<31396> A_IWL<31395> A_IWL<31394> A_IWL<31393> A_IWL<31392> A_IWL<31391> A_IWL<31390> A_IWL<31389> A_IWL<31388> A_IWL<31387> A_IWL<31386> A_IWL<31385> A_IWL<31384> A_IWL<31383> A_IWL<31382> A_IWL<31381> A_IWL<31380> A_IWL<31379> A_IWL<31378> A_IWL<31377> A_IWL<31376> A_IWL<31375> A_IWL<31374> A_IWL<31373> A_IWL<31372> A_IWL<31371> A_IWL<31370> A_IWL<31369> A_IWL<31368> A_IWL<31367> A_IWL<31366> A_IWL<31365> A_IWL<31364> A_IWL<31363> A_IWL<31362> A_IWL<31361> A_IWL<31360> A_IWL<31359> A_IWL<31358> A_IWL<31357> A_IWL<31356> A_IWL<31355> A_IWL<31354> A_IWL<31353> A_IWL<31352> A_IWL<31351> A_IWL<31350> A_IWL<31349> A_IWL<31348> A_IWL<31347> A_IWL<31346> A_IWL<31345> A_IWL<31344> A_IWL<31343> A_IWL<31342> A_IWL<31341> A_IWL<31340> A_IWL<31339> A_IWL<31338> A_IWL<31337> A_IWL<31336> A_IWL<31335> A_IWL<31334> A_IWL<31333> A_IWL<31332> A_IWL<31331> A_IWL<31330> A_IWL<31329> A_IWL<31328> A_IWL<31327> A_IWL<31326> A_IWL<31325> A_IWL<31324> A_IWL<31323> A_IWL<31322> A_IWL<31321> A_IWL<31320> A_IWL<31319> A_IWL<31318> A_IWL<31317> A_IWL<31316> A_IWL<31315> A_IWL<31314> A_IWL<31313> A_IWL<31312> A_IWL<31311> A_IWL<31310> A_IWL<31309> A_IWL<31308> A_IWL<31307> A_IWL<31306> A_IWL<31305> A_IWL<31304> A_IWL<31303> A_IWL<31302> A_IWL<31301> A_IWL<31300> A_IWL<31299> A_IWL<31298> A_IWL<31297> A_IWL<31296> A_IWL<31295> A_IWL<31294> A_IWL<31293> A_IWL<31292> A_IWL<31291> A_IWL<31290> A_IWL<31289> A_IWL<31288> A_IWL<31287> A_IWL<31286> A_IWL<31285> A_IWL<31284> A_IWL<31283> A_IWL<31282> A_IWL<31281> A_IWL<31280> A_IWL<31279> A_IWL<31278> A_IWL<31277> A_IWL<31276> A_IWL<31275> A_IWL<31274> A_IWL<31273> A_IWL<31272> A_IWL<31271> A_IWL<31270> A_IWL<31269> A_IWL<31268> A_IWL<31267> A_IWL<31266> A_IWL<31265> A_IWL<31264> A_IWL<31263> A_IWL<31262> A_IWL<31261> A_IWL<31260> A_IWL<31259> A_IWL<31258> A_IWL<31257> A_IWL<31256> A_IWL<31255> A_IWL<31254> A_IWL<31253> A_IWL<31252> A_IWL<31251> A_IWL<31250> A_IWL<31249> A_IWL<31248> A_IWL<31247> A_IWL<31246> A_IWL<31245> A_IWL<31244> A_IWL<31243> A_IWL<31242> A_IWL<31241> A_IWL<31240> A_IWL<31239> A_IWL<31238> A_IWL<31237> A_IWL<31236> A_IWL<31235> A_IWL<31234> A_IWL<31233> A_IWL<31232> A_IWL<32255> A_IWL<32254> A_IWL<32253> A_IWL<32252> A_IWL<32251> A_IWL<32250> A_IWL<32249> A_IWL<32248> A_IWL<32247> A_IWL<32246> A_IWL<32245> A_IWL<32244> A_IWL<32243> A_IWL<32242> A_IWL<32241> A_IWL<32240> A_IWL<32239> A_IWL<32238> A_IWL<32237> A_IWL<32236> A_IWL<32235> A_IWL<32234> A_IWL<32233> A_IWL<32232> A_IWL<32231> A_IWL<32230> A_IWL<32229> A_IWL<32228> A_IWL<32227> A_IWL<32226> A_IWL<32225> A_IWL<32224> A_IWL<32223> A_IWL<32222> A_IWL<32221> A_IWL<32220> A_IWL<32219> A_IWL<32218> A_IWL<32217> A_IWL<32216> A_IWL<32215> A_IWL<32214> A_IWL<32213> A_IWL<32212> A_IWL<32211> A_IWL<32210> A_IWL<32209> A_IWL<32208> A_IWL<32207> A_IWL<32206> A_IWL<32205> A_IWL<32204> A_IWL<32203> A_IWL<32202> A_IWL<32201> A_IWL<32200> A_IWL<32199> A_IWL<32198> A_IWL<32197> A_IWL<32196> A_IWL<32195> A_IWL<32194> A_IWL<32193> A_IWL<32192> A_IWL<32191> A_IWL<32190> A_IWL<32189> A_IWL<32188> A_IWL<32187> A_IWL<32186> A_IWL<32185> A_IWL<32184> A_IWL<32183> A_IWL<32182> A_IWL<32181> A_IWL<32180> A_IWL<32179> A_IWL<32178> A_IWL<32177> A_IWL<32176> A_IWL<32175> A_IWL<32174> A_IWL<32173> A_IWL<32172> A_IWL<32171> A_IWL<32170> A_IWL<32169> A_IWL<32168> A_IWL<32167> A_IWL<32166> A_IWL<32165> A_IWL<32164> A_IWL<32163> A_IWL<32162> A_IWL<32161> A_IWL<32160> A_IWL<32159> A_IWL<32158> A_IWL<32157> A_IWL<32156> A_IWL<32155> A_IWL<32154> A_IWL<32153> A_IWL<32152> A_IWL<32151> A_IWL<32150> A_IWL<32149> A_IWL<32148> A_IWL<32147> A_IWL<32146> A_IWL<32145> A_IWL<32144> A_IWL<32143> A_IWL<32142> A_IWL<32141> A_IWL<32140> A_IWL<32139> A_IWL<32138> A_IWL<32137> A_IWL<32136> A_IWL<32135> A_IWL<32134> A_IWL<32133> A_IWL<32132> A_IWL<32131> A_IWL<32130> A_IWL<32129> A_IWL<32128> A_IWL<32127> A_IWL<32126> A_IWL<32125> A_IWL<32124> A_IWL<32123> A_IWL<32122> A_IWL<32121> A_IWL<32120> A_IWL<32119> A_IWL<32118> A_IWL<32117> A_IWL<32116> A_IWL<32115> A_IWL<32114> A_IWL<32113> A_IWL<32112> A_IWL<32111> A_IWL<32110> A_IWL<32109> A_IWL<32108> A_IWL<32107> A_IWL<32106> A_IWL<32105> A_IWL<32104> A_IWL<32103> A_IWL<32102> A_IWL<32101> A_IWL<32100> A_IWL<32099> A_IWL<32098> A_IWL<32097> A_IWL<32096> A_IWL<32095> A_IWL<32094> A_IWL<32093> A_IWL<32092> A_IWL<32091> A_IWL<32090> A_IWL<32089> A_IWL<32088> A_IWL<32087> A_IWL<32086> A_IWL<32085> A_IWL<32084> A_IWL<32083> A_IWL<32082> A_IWL<32081> A_IWL<32080> A_IWL<32079> A_IWL<32078> A_IWL<32077> A_IWL<32076> A_IWL<32075> A_IWL<32074> A_IWL<32073> A_IWL<32072> A_IWL<32071> A_IWL<32070> A_IWL<32069> A_IWL<32068> A_IWL<32067> A_IWL<32066> A_IWL<32065> A_IWL<32064> A_IWL<32063> A_IWL<32062> A_IWL<32061> A_IWL<32060> A_IWL<32059> A_IWL<32058> A_IWL<32057> A_IWL<32056> A_IWL<32055> A_IWL<32054> A_IWL<32053> A_IWL<32052> A_IWL<32051> A_IWL<32050> A_IWL<32049> A_IWL<32048> A_IWL<32047> A_IWL<32046> A_IWL<32045> A_IWL<32044> A_IWL<32043> A_IWL<32042> A_IWL<32041> A_IWL<32040> A_IWL<32039> A_IWL<32038> A_IWL<32037> A_IWL<32036> A_IWL<32035> A_IWL<32034> A_IWL<32033> A_IWL<32032> A_IWL<32031> A_IWL<32030> A_IWL<32029> A_IWL<32028> A_IWL<32027> A_IWL<32026> A_IWL<32025> A_IWL<32024> A_IWL<32023> A_IWL<32022> A_IWL<32021> A_IWL<32020> A_IWL<32019> A_IWL<32018> A_IWL<32017> A_IWL<32016> A_IWL<32015> A_IWL<32014> A_IWL<32013> A_IWL<32012> A_IWL<32011> A_IWL<32010> A_IWL<32009> A_IWL<32008> A_IWL<32007> A_IWL<32006> A_IWL<32005> A_IWL<32004> A_IWL<32003> A_IWL<32002> A_IWL<32001> A_IWL<32000> A_IWL<31999> A_IWL<31998> A_IWL<31997> A_IWL<31996> A_IWL<31995> A_IWL<31994> A_IWL<31993> A_IWL<31992> A_IWL<31991> A_IWL<31990> A_IWL<31989> A_IWL<31988> A_IWL<31987> A_IWL<31986> A_IWL<31985> A_IWL<31984> A_IWL<31983> A_IWL<31982> A_IWL<31981> A_IWL<31980> A_IWL<31979> A_IWL<31978> A_IWL<31977> A_IWL<31976> A_IWL<31975> A_IWL<31974> A_IWL<31973> A_IWL<31972> A_IWL<31971> A_IWL<31970> A_IWL<31969> A_IWL<31968> A_IWL<31967> A_IWL<31966> A_IWL<31965> A_IWL<31964> A_IWL<31963> A_IWL<31962> A_IWL<31961> A_IWL<31960> A_IWL<31959> A_IWL<31958> A_IWL<31957> A_IWL<31956> A_IWL<31955> A_IWL<31954> A_IWL<31953> A_IWL<31952> A_IWL<31951> A_IWL<31950> A_IWL<31949> A_IWL<31948> A_IWL<31947> A_IWL<31946> A_IWL<31945> A_IWL<31944> A_IWL<31943> A_IWL<31942> A_IWL<31941> A_IWL<31940> A_IWL<31939> A_IWL<31938> A_IWL<31937> A_IWL<31936> A_IWL<31935> A_IWL<31934> A_IWL<31933> A_IWL<31932> A_IWL<31931> A_IWL<31930> A_IWL<31929> A_IWL<31928> A_IWL<31927> A_IWL<31926> A_IWL<31925> A_IWL<31924> A_IWL<31923> A_IWL<31922> A_IWL<31921> A_IWL<31920> A_IWL<31919> A_IWL<31918> A_IWL<31917> A_IWL<31916> A_IWL<31915> A_IWL<31914> A_IWL<31913> A_IWL<31912> A_IWL<31911> A_IWL<31910> A_IWL<31909> A_IWL<31908> A_IWL<31907> A_IWL<31906> A_IWL<31905> A_IWL<31904> A_IWL<31903> A_IWL<31902> A_IWL<31901> A_IWL<31900> A_IWL<31899> A_IWL<31898> A_IWL<31897> A_IWL<31896> A_IWL<31895> A_IWL<31894> A_IWL<31893> A_IWL<31892> A_IWL<31891> A_IWL<31890> A_IWL<31889> A_IWL<31888> A_IWL<31887> A_IWL<31886> A_IWL<31885> A_IWL<31884> A_IWL<31883> A_IWL<31882> A_IWL<31881> A_IWL<31880> A_IWL<31879> A_IWL<31878> A_IWL<31877> A_IWL<31876> A_IWL<31875> A_IWL<31874> A_IWL<31873> A_IWL<31872> A_IWL<31871> A_IWL<31870> A_IWL<31869> A_IWL<31868> A_IWL<31867> A_IWL<31866> A_IWL<31865> A_IWL<31864> A_IWL<31863> A_IWL<31862> A_IWL<31861> A_IWL<31860> A_IWL<31859> A_IWL<31858> A_IWL<31857> A_IWL<31856> A_IWL<31855> A_IWL<31854> A_IWL<31853> A_IWL<31852> A_IWL<31851> A_IWL<31850> A_IWL<31849> A_IWL<31848> A_IWL<31847> A_IWL<31846> A_IWL<31845> A_IWL<31844> A_IWL<31843> A_IWL<31842> A_IWL<31841> A_IWL<31840> A_IWL<31839> A_IWL<31838> A_IWL<31837> A_IWL<31836> A_IWL<31835> A_IWL<31834> A_IWL<31833> A_IWL<31832> A_IWL<31831> A_IWL<31830> A_IWL<31829> A_IWL<31828> A_IWL<31827> A_IWL<31826> A_IWL<31825> A_IWL<31824> A_IWL<31823> A_IWL<31822> A_IWL<31821> A_IWL<31820> A_IWL<31819> A_IWL<31818> A_IWL<31817> A_IWL<31816> A_IWL<31815> A_IWL<31814> A_IWL<31813> A_IWL<31812> A_IWL<31811> A_IWL<31810> A_IWL<31809> A_IWL<31808> A_IWL<31807> A_IWL<31806> A_IWL<31805> A_IWL<31804> A_IWL<31803> A_IWL<31802> A_IWL<31801> A_IWL<31800> A_IWL<31799> A_IWL<31798> A_IWL<31797> A_IWL<31796> A_IWL<31795> A_IWL<31794> A_IWL<31793> A_IWL<31792> A_IWL<31791> A_IWL<31790> A_IWL<31789> A_IWL<31788> A_IWL<31787> A_IWL<31786> A_IWL<31785> A_IWL<31784> A_IWL<31783> A_IWL<31782> A_IWL<31781> A_IWL<31780> A_IWL<31779> A_IWL<31778> A_IWL<31777> A_IWL<31776> A_IWL<31775> A_IWL<31774> A_IWL<31773> A_IWL<31772> A_IWL<31771> A_IWL<31770> A_IWL<31769> A_IWL<31768> A_IWL<31767> A_IWL<31766> A_IWL<31765> A_IWL<31764> A_IWL<31763> A_IWL<31762> A_IWL<31761> A_IWL<31760> A_IWL<31759> A_IWL<31758> A_IWL<31757> A_IWL<31756> A_IWL<31755> A_IWL<31754> A_IWL<31753> A_IWL<31752> A_IWL<31751> A_IWL<31750> A_IWL<31749> A_IWL<31748> A_IWL<31747> A_IWL<31746> A_IWL<31745> A_IWL<31744> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<61> A_BLC<123> A_BLC<122> A_BLC_TOP<123> A_BLC_TOP<122> A_BLT<123> A_BLT<122> A_BLT_TOP<123> A_BLT_TOP<122> A_IWL<31231> A_IWL<31230> A_IWL<31229> A_IWL<31228> A_IWL<31227> A_IWL<31226> A_IWL<31225> A_IWL<31224> A_IWL<31223> A_IWL<31222> A_IWL<31221> A_IWL<31220> A_IWL<31219> A_IWL<31218> A_IWL<31217> A_IWL<31216> A_IWL<31215> A_IWL<31214> A_IWL<31213> A_IWL<31212> A_IWL<31211> A_IWL<31210> A_IWL<31209> A_IWL<31208> A_IWL<31207> A_IWL<31206> A_IWL<31205> A_IWL<31204> A_IWL<31203> A_IWL<31202> A_IWL<31201> A_IWL<31200> A_IWL<31199> A_IWL<31198> A_IWL<31197> A_IWL<31196> A_IWL<31195> A_IWL<31194> A_IWL<31193> A_IWL<31192> A_IWL<31191> A_IWL<31190> A_IWL<31189> A_IWL<31188> A_IWL<31187> A_IWL<31186> A_IWL<31185> A_IWL<31184> A_IWL<31183> A_IWL<31182> A_IWL<31181> A_IWL<31180> A_IWL<31179> A_IWL<31178> A_IWL<31177> A_IWL<31176> A_IWL<31175> A_IWL<31174> A_IWL<31173> A_IWL<31172> A_IWL<31171> A_IWL<31170> A_IWL<31169> A_IWL<31168> A_IWL<31167> A_IWL<31166> A_IWL<31165> A_IWL<31164> A_IWL<31163> A_IWL<31162> A_IWL<31161> A_IWL<31160> A_IWL<31159> A_IWL<31158> A_IWL<31157> A_IWL<31156> A_IWL<31155> A_IWL<31154> A_IWL<31153> A_IWL<31152> A_IWL<31151> A_IWL<31150> A_IWL<31149> A_IWL<31148> A_IWL<31147> A_IWL<31146> A_IWL<31145> A_IWL<31144> A_IWL<31143> A_IWL<31142> A_IWL<31141> A_IWL<31140> A_IWL<31139> A_IWL<31138> A_IWL<31137> A_IWL<31136> A_IWL<31135> A_IWL<31134> A_IWL<31133> A_IWL<31132> A_IWL<31131> A_IWL<31130> A_IWL<31129> A_IWL<31128> A_IWL<31127> A_IWL<31126> A_IWL<31125> A_IWL<31124> A_IWL<31123> A_IWL<31122> A_IWL<31121> A_IWL<31120> A_IWL<31119> A_IWL<31118> A_IWL<31117> A_IWL<31116> A_IWL<31115> A_IWL<31114> A_IWL<31113> A_IWL<31112> A_IWL<31111> A_IWL<31110> A_IWL<31109> A_IWL<31108> A_IWL<31107> A_IWL<31106> A_IWL<31105> A_IWL<31104> A_IWL<31103> A_IWL<31102> A_IWL<31101> A_IWL<31100> A_IWL<31099> A_IWL<31098> A_IWL<31097> A_IWL<31096> A_IWL<31095> A_IWL<31094> A_IWL<31093> A_IWL<31092> A_IWL<31091> A_IWL<31090> A_IWL<31089> A_IWL<31088> A_IWL<31087> A_IWL<31086> A_IWL<31085> A_IWL<31084> A_IWL<31083> A_IWL<31082> A_IWL<31081> A_IWL<31080> A_IWL<31079> A_IWL<31078> A_IWL<31077> A_IWL<31076> A_IWL<31075> A_IWL<31074> A_IWL<31073> A_IWL<31072> A_IWL<31071> A_IWL<31070> A_IWL<31069> A_IWL<31068> A_IWL<31067> A_IWL<31066> A_IWL<31065> A_IWL<31064> A_IWL<31063> A_IWL<31062> A_IWL<31061> A_IWL<31060> A_IWL<31059> A_IWL<31058> A_IWL<31057> A_IWL<31056> A_IWL<31055> A_IWL<31054> A_IWL<31053> A_IWL<31052> A_IWL<31051> A_IWL<31050> A_IWL<31049> A_IWL<31048> A_IWL<31047> A_IWL<31046> A_IWL<31045> A_IWL<31044> A_IWL<31043> A_IWL<31042> A_IWL<31041> A_IWL<31040> A_IWL<31039> A_IWL<31038> A_IWL<31037> A_IWL<31036> A_IWL<31035> A_IWL<31034> A_IWL<31033> A_IWL<31032> A_IWL<31031> A_IWL<31030> A_IWL<31029> A_IWL<31028> A_IWL<31027> A_IWL<31026> A_IWL<31025> A_IWL<31024> A_IWL<31023> A_IWL<31022> A_IWL<31021> A_IWL<31020> A_IWL<31019> A_IWL<31018> A_IWL<31017> A_IWL<31016> A_IWL<31015> A_IWL<31014> A_IWL<31013> A_IWL<31012> A_IWL<31011> A_IWL<31010> A_IWL<31009> A_IWL<31008> A_IWL<31007> A_IWL<31006> A_IWL<31005> A_IWL<31004> A_IWL<31003> A_IWL<31002> A_IWL<31001> A_IWL<31000> A_IWL<30999> A_IWL<30998> A_IWL<30997> A_IWL<30996> A_IWL<30995> A_IWL<30994> A_IWL<30993> A_IWL<30992> A_IWL<30991> A_IWL<30990> A_IWL<30989> A_IWL<30988> A_IWL<30987> A_IWL<30986> A_IWL<30985> A_IWL<30984> A_IWL<30983> A_IWL<30982> A_IWL<30981> A_IWL<30980> A_IWL<30979> A_IWL<30978> A_IWL<30977> A_IWL<30976> A_IWL<30975> A_IWL<30974> A_IWL<30973> A_IWL<30972> A_IWL<30971> A_IWL<30970> A_IWL<30969> A_IWL<30968> A_IWL<30967> A_IWL<30966> A_IWL<30965> A_IWL<30964> A_IWL<30963> A_IWL<30962> A_IWL<30961> A_IWL<30960> A_IWL<30959> A_IWL<30958> A_IWL<30957> A_IWL<30956> A_IWL<30955> A_IWL<30954> A_IWL<30953> A_IWL<30952> A_IWL<30951> A_IWL<30950> A_IWL<30949> A_IWL<30948> A_IWL<30947> A_IWL<30946> A_IWL<30945> A_IWL<30944> A_IWL<30943> A_IWL<30942> A_IWL<30941> A_IWL<30940> A_IWL<30939> A_IWL<30938> A_IWL<30937> A_IWL<30936> A_IWL<30935> A_IWL<30934> A_IWL<30933> A_IWL<30932> A_IWL<30931> A_IWL<30930> A_IWL<30929> A_IWL<30928> A_IWL<30927> A_IWL<30926> A_IWL<30925> A_IWL<30924> A_IWL<30923> A_IWL<30922> A_IWL<30921> A_IWL<30920> A_IWL<30919> A_IWL<30918> A_IWL<30917> A_IWL<30916> A_IWL<30915> A_IWL<30914> A_IWL<30913> A_IWL<30912> A_IWL<30911> A_IWL<30910> A_IWL<30909> A_IWL<30908> A_IWL<30907> A_IWL<30906> A_IWL<30905> A_IWL<30904> A_IWL<30903> A_IWL<30902> A_IWL<30901> A_IWL<30900> A_IWL<30899> A_IWL<30898> A_IWL<30897> A_IWL<30896> A_IWL<30895> A_IWL<30894> A_IWL<30893> A_IWL<30892> A_IWL<30891> A_IWL<30890> A_IWL<30889> A_IWL<30888> A_IWL<30887> A_IWL<30886> A_IWL<30885> A_IWL<30884> A_IWL<30883> A_IWL<30882> A_IWL<30881> A_IWL<30880> A_IWL<30879> A_IWL<30878> A_IWL<30877> A_IWL<30876> A_IWL<30875> A_IWL<30874> A_IWL<30873> A_IWL<30872> A_IWL<30871> A_IWL<30870> A_IWL<30869> A_IWL<30868> A_IWL<30867> A_IWL<30866> A_IWL<30865> A_IWL<30864> A_IWL<30863> A_IWL<30862> A_IWL<30861> A_IWL<30860> A_IWL<30859> A_IWL<30858> A_IWL<30857> A_IWL<30856> A_IWL<30855> A_IWL<30854> A_IWL<30853> A_IWL<30852> A_IWL<30851> A_IWL<30850> A_IWL<30849> A_IWL<30848> A_IWL<30847> A_IWL<30846> A_IWL<30845> A_IWL<30844> A_IWL<30843> A_IWL<30842> A_IWL<30841> A_IWL<30840> A_IWL<30839> A_IWL<30838> A_IWL<30837> A_IWL<30836> A_IWL<30835> A_IWL<30834> A_IWL<30833> A_IWL<30832> A_IWL<30831> A_IWL<30830> A_IWL<30829> A_IWL<30828> A_IWL<30827> A_IWL<30826> A_IWL<30825> A_IWL<30824> A_IWL<30823> A_IWL<30822> A_IWL<30821> A_IWL<30820> A_IWL<30819> A_IWL<30818> A_IWL<30817> A_IWL<30816> A_IWL<30815> A_IWL<30814> A_IWL<30813> A_IWL<30812> A_IWL<30811> A_IWL<30810> A_IWL<30809> A_IWL<30808> A_IWL<30807> A_IWL<30806> A_IWL<30805> A_IWL<30804> A_IWL<30803> A_IWL<30802> A_IWL<30801> A_IWL<30800> A_IWL<30799> A_IWL<30798> A_IWL<30797> A_IWL<30796> A_IWL<30795> A_IWL<30794> A_IWL<30793> A_IWL<30792> A_IWL<30791> A_IWL<30790> A_IWL<30789> A_IWL<30788> A_IWL<30787> A_IWL<30786> A_IWL<30785> A_IWL<30784> A_IWL<30783> A_IWL<30782> A_IWL<30781> A_IWL<30780> A_IWL<30779> A_IWL<30778> A_IWL<30777> A_IWL<30776> A_IWL<30775> A_IWL<30774> A_IWL<30773> A_IWL<30772> A_IWL<30771> A_IWL<30770> A_IWL<30769> A_IWL<30768> A_IWL<30767> A_IWL<30766> A_IWL<30765> A_IWL<30764> A_IWL<30763> A_IWL<30762> A_IWL<30761> A_IWL<30760> A_IWL<30759> A_IWL<30758> A_IWL<30757> A_IWL<30756> A_IWL<30755> A_IWL<30754> A_IWL<30753> A_IWL<30752> A_IWL<30751> A_IWL<30750> A_IWL<30749> A_IWL<30748> A_IWL<30747> A_IWL<30746> A_IWL<30745> A_IWL<30744> A_IWL<30743> A_IWL<30742> A_IWL<30741> A_IWL<30740> A_IWL<30739> A_IWL<30738> A_IWL<30737> A_IWL<30736> A_IWL<30735> A_IWL<30734> A_IWL<30733> A_IWL<30732> A_IWL<30731> A_IWL<30730> A_IWL<30729> A_IWL<30728> A_IWL<30727> A_IWL<30726> A_IWL<30725> A_IWL<30724> A_IWL<30723> A_IWL<30722> A_IWL<30721> A_IWL<30720> A_IWL<31743> A_IWL<31742> A_IWL<31741> A_IWL<31740> A_IWL<31739> A_IWL<31738> A_IWL<31737> A_IWL<31736> A_IWL<31735> A_IWL<31734> A_IWL<31733> A_IWL<31732> A_IWL<31731> A_IWL<31730> A_IWL<31729> A_IWL<31728> A_IWL<31727> A_IWL<31726> A_IWL<31725> A_IWL<31724> A_IWL<31723> A_IWL<31722> A_IWL<31721> A_IWL<31720> A_IWL<31719> A_IWL<31718> A_IWL<31717> A_IWL<31716> A_IWL<31715> A_IWL<31714> A_IWL<31713> A_IWL<31712> A_IWL<31711> A_IWL<31710> A_IWL<31709> A_IWL<31708> A_IWL<31707> A_IWL<31706> A_IWL<31705> A_IWL<31704> A_IWL<31703> A_IWL<31702> A_IWL<31701> A_IWL<31700> A_IWL<31699> A_IWL<31698> A_IWL<31697> A_IWL<31696> A_IWL<31695> A_IWL<31694> A_IWL<31693> A_IWL<31692> A_IWL<31691> A_IWL<31690> A_IWL<31689> A_IWL<31688> A_IWL<31687> A_IWL<31686> A_IWL<31685> A_IWL<31684> A_IWL<31683> A_IWL<31682> A_IWL<31681> A_IWL<31680> A_IWL<31679> A_IWL<31678> A_IWL<31677> A_IWL<31676> A_IWL<31675> A_IWL<31674> A_IWL<31673> A_IWL<31672> A_IWL<31671> A_IWL<31670> A_IWL<31669> A_IWL<31668> A_IWL<31667> A_IWL<31666> A_IWL<31665> A_IWL<31664> A_IWL<31663> A_IWL<31662> A_IWL<31661> A_IWL<31660> A_IWL<31659> A_IWL<31658> A_IWL<31657> A_IWL<31656> A_IWL<31655> A_IWL<31654> A_IWL<31653> A_IWL<31652> A_IWL<31651> A_IWL<31650> A_IWL<31649> A_IWL<31648> A_IWL<31647> A_IWL<31646> A_IWL<31645> A_IWL<31644> A_IWL<31643> A_IWL<31642> A_IWL<31641> A_IWL<31640> A_IWL<31639> A_IWL<31638> A_IWL<31637> A_IWL<31636> A_IWL<31635> A_IWL<31634> A_IWL<31633> A_IWL<31632> A_IWL<31631> A_IWL<31630> A_IWL<31629> A_IWL<31628> A_IWL<31627> A_IWL<31626> A_IWL<31625> A_IWL<31624> A_IWL<31623> A_IWL<31622> A_IWL<31621> A_IWL<31620> A_IWL<31619> A_IWL<31618> A_IWL<31617> A_IWL<31616> A_IWL<31615> A_IWL<31614> A_IWL<31613> A_IWL<31612> A_IWL<31611> A_IWL<31610> A_IWL<31609> A_IWL<31608> A_IWL<31607> A_IWL<31606> A_IWL<31605> A_IWL<31604> A_IWL<31603> A_IWL<31602> A_IWL<31601> A_IWL<31600> A_IWL<31599> A_IWL<31598> A_IWL<31597> A_IWL<31596> A_IWL<31595> A_IWL<31594> A_IWL<31593> A_IWL<31592> A_IWL<31591> A_IWL<31590> A_IWL<31589> A_IWL<31588> A_IWL<31587> A_IWL<31586> A_IWL<31585> A_IWL<31584> A_IWL<31583> A_IWL<31582> A_IWL<31581> A_IWL<31580> A_IWL<31579> A_IWL<31578> A_IWL<31577> A_IWL<31576> A_IWL<31575> A_IWL<31574> A_IWL<31573> A_IWL<31572> A_IWL<31571> A_IWL<31570> A_IWL<31569> A_IWL<31568> A_IWL<31567> A_IWL<31566> A_IWL<31565> A_IWL<31564> A_IWL<31563> A_IWL<31562> A_IWL<31561> A_IWL<31560> A_IWL<31559> A_IWL<31558> A_IWL<31557> A_IWL<31556> A_IWL<31555> A_IWL<31554> A_IWL<31553> A_IWL<31552> A_IWL<31551> A_IWL<31550> A_IWL<31549> A_IWL<31548> A_IWL<31547> A_IWL<31546> A_IWL<31545> A_IWL<31544> A_IWL<31543> A_IWL<31542> A_IWL<31541> A_IWL<31540> A_IWL<31539> A_IWL<31538> A_IWL<31537> A_IWL<31536> A_IWL<31535> A_IWL<31534> A_IWL<31533> A_IWL<31532> A_IWL<31531> A_IWL<31530> A_IWL<31529> A_IWL<31528> A_IWL<31527> A_IWL<31526> A_IWL<31525> A_IWL<31524> A_IWL<31523> A_IWL<31522> A_IWL<31521> A_IWL<31520> A_IWL<31519> A_IWL<31518> A_IWL<31517> A_IWL<31516> A_IWL<31515> A_IWL<31514> A_IWL<31513> A_IWL<31512> A_IWL<31511> A_IWL<31510> A_IWL<31509> A_IWL<31508> A_IWL<31507> A_IWL<31506> A_IWL<31505> A_IWL<31504> A_IWL<31503> A_IWL<31502> A_IWL<31501> A_IWL<31500> A_IWL<31499> A_IWL<31498> A_IWL<31497> A_IWL<31496> A_IWL<31495> A_IWL<31494> A_IWL<31493> A_IWL<31492> A_IWL<31491> A_IWL<31490> A_IWL<31489> A_IWL<31488> A_IWL<31487> A_IWL<31486> A_IWL<31485> A_IWL<31484> A_IWL<31483> A_IWL<31482> A_IWL<31481> A_IWL<31480> A_IWL<31479> A_IWL<31478> A_IWL<31477> A_IWL<31476> A_IWL<31475> A_IWL<31474> A_IWL<31473> A_IWL<31472> A_IWL<31471> A_IWL<31470> A_IWL<31469> A_IWL<31468> A_IWL<31467> A_IWL<31466> A_IWL<31465> A_IWL<31464> A_IWL<31463> A_IWL<31462> A_IWL<31461> A_IWL<31460> A_IWL<31459> A_IWL<31458> A_IWL<31457> A_IWL<31456> A_IWL<31455> A_IWL<31454> A_IWL<31453> A_IWL<31452> A_IWL<31451> A_IWL<31450> A_IWL<31449> A_IWL<31448> A_IWL<31447> A_IWL<31446> A_IWL<31445> A_IWL<31444> A_IWL<31443> A_IWL<31442> A_IWL<31441> A_IWL<31440> A_IWL<31439> A_IWL<31438> A_IWL<31437> A_IWL<31436> A_IWL<31435> A_IWL<31434> A_IWL<31433> A_IWL<31432> A_IWL<31431> A_IWL<31430> A_IWL<31429> A_IWL<31428> A_IWL<31427> A_IWL<31426> A_IWL<31425> A_IWL<31424> A_IWL<31423> A_IWL<31422> A_IWL<31421> A_IWL<31420> A_IWL<31419> A_IWL<31418> A_IWL<31417> A_IWL<31416> A_IWL<31415> A_IWL<31414> A_IWL<31413> A_IWL<31412> A_IWL<31411> A_IWL<31410> A_IWL<31409> A_IWL<31408> A_IWL<31407> A_IWL<31406> A_IWL<31405> A_IWL<31404> A_IWL<31403> A_IWL<31402> A_IWL<31401> A_IWL<31400> A_IWL<31399> A_IWL<31398> A_IWL<31397> A_IWL<31396> A_IWL<31395> A_IWL<31394> A_IWL<31393> A_IWL<31392> A_IWL<31391> A_IWL<31390> A_IWL<31389> A_IWL<31388> A_IWL<31387> A_IWL<31386> A_IWL<31385> A_IWL<31384> A_IWL<31383> A_IWL<31382> A_IWL<31381> A_IWL<31380> A_IWL<31379> A_IWL<31378> A_IWL<31377> A_IWL<31376> A_IWL<31375> A_IWL<31374> A_IWL<31373> A_IWL<31372> A_IWL<31371> A_IWL<31370> A_IWL<31369> A_IWL<31368> A_IWL<31367> A_IWL<31366> A_IWL<31365> A_IWL<31364> A_IWL<31363> A_IWL<31362> A_IWL<31361> A_IWL<31360> A_IWL<31359> A_IWL<31358> A_IWL<31357> A_IWL<31356> A_IWL<31355> A_IWL<31354> A_IWL<31353> A_IWL<31352> A_IWL<31351> A_IWL<31350> A_IWL<31349> A_IWL<31348> A_IWL<31347> A_IWL<31346> A_IWL<31345> A_IWL<31344> A_IWL<31343> A_IWL<31342> A_IWL<31341> A_IWL<31340> A_IWL<31339> A_IWL<31338> A_IWL<31337> A_IWL<31336> A_IWL<31335> A_IWL<31334> A_IWL<31333> A_IWL<31332> A_IWL<31331> A_IWL<31330> A_IWL<31329> A_IWL<31328> A_IWL<31327> A_IWL<31326> A_IWL<31325> A_IWL<31324> A_IWL<31323> A_IWL<31322> A_IWL<31321> A_IWL<31320> A_IWL<31319> A_IWL<31318> A_IWL<31317> A_IWL<31316> A_IWL<31315> A_IWL<31314> A_IWL<31313> A_IWL<31312> A_IWL<31311> A_IWL<31310> A_IWL<31309> A_IWL<31308> A_IWL<31307> A_IWL<31306> A_IWL<31305> A_IWL<31304> A_IWL<31303> A_IWL<31302> A_IWL<31301> A_IWL<31300> A_IWL<31299> A_IWL<31298> A_IWL<31297> A_IWL<31296> A_IWL<31295> A_IWL<31294> A_IWL<31293> A_IWL<31292> A_IWL<31291> A_IWL<31290> A_IWL<31289> A_IWL<31288> A_IWL<31287> A_IWL<31286> A_IWL<31285> A_IWL<31284> A_IWL<31283> A_IWL<31282> A_IWL<31281> A_IWL<31280> A_IWL<31279> A_IWL<31278> A_IWL<31277> A_IWL<31276> A_IWL<31275> A_IWL<31274> A_IWL<31273> A_IWL<31272> A_IWL<31271> A_IWL<31270> A_IWL<31269> A_IWL<31268> A_IWL<31267> A_IWL<31266> A_IWL<31265> A_IWL<31264> A_IWL<31263> A_IWL<31262> A_IWL<31261> A_IWL<31260> A_IWL<31259> A_IWL<31258> A_IWL<31257> A_IWL<31256> A_IWL<31255> A_IWL<31254> A_IWL<31253> A_IWL<31252> A_IWL<31251> A_IWL<31250> A_IWL<31249> A_IWL<31248> A_IWL<31247> A_IWL<31246> A_IWL<31245> A_IWL<31244> A_IWL<31243> A_IWL<31242> A_IWL<31241> A_IWL<31240> A_IWL<31239> A_IWL<31238> A_IWL<31237> A_IWL<31236> A_IWL<31235> A_IWL<31234> A_IWL<31233> A_IWL<31232> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<60> A_BLC<121> A_BLC<120> A_BLC_TOP<121> A_BLC_TOP<120> A_BLT<121> A_BLT<120> A_BLT_TOP<121> A_BLT_TOP<120> A_IWL<30719> A_IWL<30718> A_IWL<30717> A_IWL<30716> A_IWL<30715> A_IWL<30714> A_IWL<30713> A_IWL<30712> A_IWL<30711> A_IWL<30710> A_IWL<30709> A_IWL<30708> A_IWL<30707> A_IWL<30706> A_IWL<30705> A_IWL<30704> A_IWL<30703> A_IWL<30702> A_IWL<30701> A_IWL<30700> A_IWL<30699> A_IWL<30698> A_IWL<30697> A_IWL<30696> A_IWL<30695> A_IWL<30694> A_IWL<30693> A_IWL<30692> A_IWL<30691> A_IWL<30690> A_IWL<30689> A_IWL<30688> A_IWL<30687> A_IWL<30686> A_IWL<30685> A_IWL<30684> A_IWL<30683> A_IWL<30682> A_IWL<30681> A_IWL<30680> A_IWL<30679> A_IWL<30678> A_IWL<30677> A_IWL<30676> A_IWL<30675> A_IWL<30674> A_IWL<30673> A_IWL<30672> A_IWL<30671> A_IWL<30670> A_IWL<30669> A_IWL<30668> A_IWL<30667> A_IWL<30666> A_IWL<30665> A_IWL<30664> A_IWL<30663> A_IWL<30662> A_IWL<30661> A_IWL<30660> A_IWL<30659> A_IWL<30658> A_IWL<30657> A_IWL<30656> A_IWL<30655> A_IWL<30654> A_IWL<30653> A_IWL<30652> A_IWL<30651> A_IWL<30650> A_IWL<30649> A_IWL<30648> A_IWL<30647> A_IWL<30646> A_IWL<30645> A_IWL<30644> A_IWL<30643> A_IWL<30642> A_IWL<30641> A_IWL<30640> A_IWL<30639> A_IWL<30638> A_IWL<30637> A_IWL<30636> A_IWL<30635> A_IWL<30634> A_IWL<30633> A_IWL<30632> A_IWL<30631> A_IWL<30630> A_IWL<30629> A_IWL<30628> A_IWL<30627> A_IWL<30626> A_IWL<30625> A_IWL<30624> A_IWL<30623> A_IWL<30622> A_IWL<30621> A_IWL<30620> A_IWL<30619> A_IWL<30618> A_IWL<30617> A_IWL<30616> A_IWL<30615> A_IWL<30614> A_IWL<30613> A_IWL<30612> A_IWL<30611> A_IWL<30610> A_IWL<30609> A_IWL<30608> A_IWL<30607> A_IWL<30606> A_IWL<30605> A_IWL<30604> A_IWL<30603> A_IWL<30602> A_IWL<30601> A_IWL<30600> A_IWL<30599> A_IWL<30598> A_IWL<30597> A_IWL<30596> A_IWL<30595> A_IWL<30594> A_IWL<30593> A_IWL<30592> A_IWL<30591> A_IWL<30590> A_IWL<30589> A_IWL<30588> A_IWL<30587> A_IWL<30586> A_IWL<30585> A_IWL<30584> A_IWL<30583> A_IWL<30582> A_IWL<30581> A_IWL<30580> A_IWL<30579> A_IWL<30578> A_IWL<30577> A_IWL<30576> A_IWL<30575> A_IWL<30574> A_IWL<30573> A_IWL<30572> A_IWL<30571> A_IWL<30570> A_IWL<30569> A_IWL<30568> A_IWL<30567> A_IWL<30566> A_IWL<30565> A_IWL<30564> A_IWL<30563> A_IWL<30562> A_IWL<30561> A_IWL<30560> A_IWL<30559> A_IWL<30558> A_IWL<30557> A_IWL<30556> A_IWL<30555> A_IWL<30554> A_IWL<30553> A_IWL<30552> A_IWL<30551> A_IWL<30550> A_IWL<30549> A_IWL<30548> A_IWL<30547> A_IWL<30546> A_IWL<30545> A_IWL<30544> A_IWL<30543> A_IWL<30542> A_IWL<30541> A_IWL<30540> A_IWL<30539> A_IWL<30538> A_IWL<30537> A_IWL<30536> A_IWL<30535> A_IWL<30534> A_IWL<30533> A_IWL<30532> A_IWL<30531> A_IWL<30530> A_IWL<30529> A_IWL<30528> A_IWL<30527> A_IWL<30526> A_IWL<30525> A_IWL<30524> A_IWL<30523> A_IWL<30522> A_IWL<30521> A_IWL<30520> A_IWL<30519> A_IWL<30518> A_IWL<30517> A_IWL<30516> A_IWL<30515> A_IWL<30514> A_IWL<30513> A_IWL<30512> A_IWL<30511> A_IWL<30510> A_IWL<30509> A_IWL<30508> A_IWL<30507> A_IWL<30506> A_IWL<30505> A_IWL<30504> A_IWL<30503> A_IWL<30502> A_IWL<30501> A_IWL<30500> A_IWL<30499> A_IWL<30498> A_IWL<30497> A_IWL<30496> A_IWL<30495> A_IWL<30494> A_IWL<30493> A_IWL<30492> A_IWL<30491> A_IWL<30490> A_IWL<30489> A_IWL<30488> A_IWL<30487> A_IWL<30486> A_IWL<30485> A_IWL<30484> A_IWL<30483> A_IWL<30482> A_IWL<30481> A_IWL<30480> A_IWL<30479> A_IWL<30478> A_IWL<30477> A_IWL<30476> A_IWL<30475> A_IWL<30474> A_IWL<30473> A_IWL<30472> A_IWL<30471> A_IWL<30470> A_IWL<30469> A_IWL<30468> A_IWL<30467> A_IWL<30466> A_IWL<30465> A_IWL<30464> A_IWL<30463> A_IWL<30462> A_IWL<30461> A_IWL<30460> A_IWL<30459> A_IWL<30458> A_IWL<30457> A_IWL<30456> A_IWL<30455> A_IWL<30454> A_IWL<30453> A_IWL<30452> A_IWL<30451> A_IWL<30450> A_IWL<30449> A_IWL<30448> A_IWL<30447> A_IWL<30446> A_IWL<30445> A_IWL<30444> A_IWL<30443> A_IWL<30442> A_IWL<30441> A_IWL<30440> A_IWL<30439> A_IWL<30438> A_IWL<30437> A_IWL<30436> A_IWL<30435> A_IWL<30434> A_IWL<30433> A_IWL<30432> A_IWL<30431> A_IWL<30430> A_IWL<30429> A_IWL<30428> A_IWL<30427> A_IWL<30426> A_IWL<30425> A_IWL<30424> A_IWL<30423> A_IWL<30422> A_IWL<30421> A_IWL<30420> A_IWL<30419> A_IWL<30418> A_IWL<30417> A_IWL<30416> A_IWL<30415> A_IWL<30414> A_IWL<30413> A_IWL<30412> A_IWL<30411> A_IWL<30410> A_IWL<30409> A_IWL<30408> A_IWL<30407> A_IWL<30406> A_IWL<30405> A_IWL<30404> A_IWL<30403> A_IWL<30402> A_IWL<30401> A_IWL<30400> A_IWL<30399> A_IWL<30398> A_IWL<30397> A_IWL<30396> A_IWL<30395> A_IWL<30394> A_IWL<30393> A_IWL<30392> A_IWL<30391> A_IWL<30390> A_IWL<30389> A_IWL<30388> A_IWL<30387> A_IWL<30386> A_IWL<30385> A_IWL<30384> A_IWL<30383> A_IWL<30382> A_IWL<30381> A_IWL<30380> A_IWL<30379> A_IWL<30378> A_IWL<30377> A_IWL<30376> A_IWL<30375> A_IWL<30374> A_IWL<30373> A_IWL<30372> A_IWL<30371> A_IWL<30370> A_IWL<30369> A_IWL<30368> A_IWL<30367> A_IWL<30366> A_IWL<30365> A_IWL<30364> A_IWL<30363> A_IWL<30362> A_IWL<30361> A_IWL<30360> A_IWL<30359> A_IWL<30358> A_IWL<30357> A_IWL<30356> A_IWL<30355> A_IWL<30354> A_IWL<30353> A_IWL<30352> A_IWL<30351> A_IWL<30350> A_IWL<30349> A_IWL<30348> A_IWL<30347> A_IWL<30346> A_IWL<30345> A_IWL<30344> A_IWL<30343> A_IWL<30342> A_IWL<30341> A_IWL<30340> A_IWL<30339> A_IWL<30338> A_IWL<30337> A_IWL<30336> A_IWL<30335> A_IWL<30334> A_IWL<30333> A_IWL<30332> A_IWL<30331> A_IWL<30330> A_IWL<30329> A_IWL<30328> A_IWL<30327> A_IWL<30326> A_IWL<30325> A_IWL<30324> A_IWL<30323> A_IWL<30322> A_IWL<30321> A_IWL<30320> A_IWL<30319> A_IWL<30318> A_IWL<30317> A_IWL<30316> A_IWL<30315> A_IWL<30314> A_IWL<30313> A_IWL<30312> A_IWL<30311> A_IWL<30310> A_IWL<30309> A_IWL<30308> A_IWL<30307> A_IWL<30306> A_IWL<30305> A_IWL<30304> A_IWL<30303> A_IWL<30302> A_IWL<30301> A_IWL<30300> A_IWL<30299> A_IWL<30298> A_IWL<30297> A_IWL<30296> A_IWL<30295> A_IWL<30294> A_IWL<30293> A_IWL<30292> A_IWL<30291> A_IWL<30290> A_IWL<30289> A_IWL<30288> A_IWL<30287> A_IWL<30286> A_IWL<30285> A_IWL<30284> A_IWL<30283> A_IWL<30282> A_IWL<30281> A_IWL<30280> A_IWL<30279> A_IWL<30278> A_IWL<30277> A_IWL<30276> A_IWL<30275> A_IWL<30274> A_IWL<30273> A_IWL<30272> A_IWL<30271> A_IWL<30270> A_IWL<30269> A_IWL<30268> A_IWL<30267> A_IWL<30266> A_IWL<30265> A_IWL<30264> A_IWL<30263> A_IWL<30262> A_IWL<30261> A_IWL<30260> A_IWL<30259> A_IWL<30258> A_IWL<30257> A_IWL<30256> A_IWL<30255> A_IWL<30254> A_IWL<30253> A_IWL<30252> A_IWL<30251> A_IWL<30250> A_IWL<30249> A_IWL<30248> A_IWL<30247> A_IWL<30246> A_IWL<30245> A_IWL<30244> A_IWL<30243> A_IWL<30242> A_IWL<30241> A_IWL<30240> A_IWL<30239> A_IWL<30238> A_IWL<30237> A_IWL<30236> A_IWL<30235> A_IWL<30234> A_IWL<30233> A_IWL<30232> A_IWL<30231> A_IWL<30230> A_IWL<30229> A_IWL<30228> A_IWL<30227> A_IWL<30226> A_IWL<30225> A_IWL<30224> A_IWL<30223> A_IWL<30222> A_IWL<30221> A_IWL<30220> A_IWL<30219> A_IWL<30218> A_IWL<30217> A_IWL<30216> A_IWL<30215> A_IWL<30214> A_IWL<30213> A_IWL<30212> A_IWL<30211> A_IWL<30210> A_IWL<30209> A_IWL<30208> A_IWL<31231> A_IWL<31230> A_IWL<31229> A_IWL<31228> A_IWL<31227> A_IWL<31226> A_IWL<31225> A_IWL<31224> A_IWL<31223> A_IWL<31222> A_IWL<31221> A_IWL<31220> A_IWL<31219> A_IWL<31218> A_IWL<31217> A_IWL<31216> A_IWL<31215> A_IWL<31214> A_IWL<31213> A_IWL<31212> A_IWL<31211> A_IWL<31210> A_IWL<31209> A_IWL<31208> A_IWL<31207> A_IWL<31206> A_IWL<31205> A_IWL<31204> A_IWL<31203> A_IWL<31202> A_IWL<31201> A_IWL<31200> A_IWL<31199> A_IWL<31198> A_IWL<31197> A_IWL<31196> A_IWL<31195> A_IWL<31194> A_IWL<31193> A_IWL<31192> A_IWL<31191> A_IWL<31190> A_IWL<31189> A_IWL<31188> A_IWL<31187> A_IWL<31186> A_IWL<31185> A_IWL<31184> A_IWL<31183> A_IWL<31182> A_IWL<31181> A_IWL<31180> A_IWL<31179> A_IWL<31178> A_IWL<31177> A_IWL<31176> A_IWL<31175> A_IWL<31174> A_IWL<31173> A_IWL<31172> A_IWL<31171> A_IWL<31170> A_IWL<31169> A_IWL<31168> A_IWL<31167> A_IWL<31166> A_IWL<31165> A_IWL<31164> A_IWL<31163> A_IWL<31162> A_IWL<31161> A_IWL<31160> A_IWL<31159> A_IWL<31158> A_IWL<31157> A_IWL<31156> A_IWL<31155> A_IWL<31154> A_IWL<31153> A_IWL<31152> A_IWL<31151> A_IWL<31150> A_IWL<31149> A_IWL<31148> A_IWL<31147> A_IWL<31146> A_IWL<31145> A_IWL<31144> A_IWL<31143> A_IWL<31142> A_IWL<31141> A_IWL<31140> A_IWL<31139> A_IWL<31138> A_IWL<31137> A_IWL<31136> A_IWL<31135> A_IWL<31134> A_IWL<31133> A_IWL<31132> A_IWL<31131> A_IWL<31130> A_IWL<31129> A_IWL<31128> A_IWL<31127> A_IWL<31126> A_IWL<31125> A_IWL<31124> A_IWL<31123> A_IWL<31122> A_IWL<31121> A_IWL<31120> A_IWL<31119> A_IWL<31118> A_IWL<31117> A_IWL<31116> A_IWL<31115> A_IWL<31114> A_IWL<31113> A_IWL<31112> A_IWL<31111> A_IWL<31110> A_IWL<31109> A_IWL<31108> A_IWL<31107> A_IWL<31106> A_IWL<31105> A_IWL<31104> A_IWL<31103> A_IWL<31102> A_IWL<31101> A_IWL<31100> A_IWL<31099> A_IWL<31098> A_IWL<31097> A_IWL<31096> A_IWL<31095> A_IWL<31094> A_IWL<31093> A_IWL<31092> A_IWL<31091> A_IWL<31090> A_IWL<31089> A_IWL<31088> A_IWL<31087> A_IWL<31086> A_IWL<31085> A_IWL<31084> A_IWL<31083> A_IWL<31082> A_IWL<31081> A_IWL<31080> A_IWL<31079> A_IWL<31078> A_IWL<31077> A_IWL<31076> A_IWL<31075> A_IWL<31074> A_IWL<31073> A_IWL<31072> A_IWL<31071> A_IWL<31070> A_IWL<31069> A_IWL<31068> A_IWL<31067> A_IWL<31066> A_IWL<31065> A_IWL<31064> A_IWL<31063> A_IWL<31062> A_IWL<31061> A_IWL<31060> A_IWL<31059> A_IWL<31058> A_IWL<31057> A_IWL<31056> A_IWL<31055> A_IWL<31054> A_IWL<31053> A_IWL<31052> A_IWL<31051> A_IWL<31050> A_IWL<31049> A_IWL<31048> A_IWL<31047> A_IWL<31046> A_IWL<31045> A_IWL<31044> A_IWL<31043> A_IWL<31042> A_IWL<31041> A_IWL<31040> A_IWL<31039> A_IWL<31038> A_IWL<31037> A_IWL<31036> A_IWL<31035> A_IWL<31034> A_IWL<31033> A_IWL<31032> A_IWL<31031> A_IWL<31030> A_IWL<31029> A_IWL<31028> A_IWL<31027> A_IWL<31026> A_IWL<31025> A_IWL<31024> A_IWL<31023> A_IWL<31022> A_IWL<31021> A_IWL<31020> A_IWL<31019> A_IWL<31018> A_IWL<31017> A_IWL<31016> A_IWL<31015> A_IWL<31014> A_IWL<31013> A_IWL<31012> A_IWL<31011> A_IWL<31010> A_IWL<31009> A_IWL<31008> A_IWL<31007> A_IWL<31006> A_IWL<31005> A_IWL<31004> A_IWL<31003> A_IWL<31002> A_IWL<31001> A_IWL<31000> A_IWL<30999> A_IWL<30998> A_IWL<30997> A_IWL<30996> A_IWL<30995> A_IWL<30994> A_IWL<30993> A_IWL<30992> A_IWL<30991> A_IWL<30990> A_IWL<30989> A_IWL<30988> A_IWL<30987> A_IWL<30986> A_IWL<30985> A_IWL<30984> A_IWL<30983> A_IWL<30982> A_IWL<30981> A_IWL<30980> A_IWL<30979> A_IWL<30978> A_IWL<30977> A_IWL<30976> A_IWL<30975> A_IWL<30974> A_IWL<30973> A_IWL<30972> A_IWL<30971> A_IWL<30970> A_IWL<30969> A_IWL<30968> A_IWL<30967> A_IWL<30966> A_IWL<30965> A_IWL<30964> A_IWL<30963> A_IWL<30962> A_IWL<30961> A_IWL<30960> A_IWL<30959> A_IWL<30958> A_IWL<30957> A_IWL<30956> A_IWL<30955> A_IWL<30954> A_IWL<30953> A_IWL<30952> A_IWL<30951> A_IWL<30950> A_IWL<30949> A_IWL<30948> A_IWL<30947> A_IWL<30946> A_IWL<30945> A_IWL<30944> A_IWL<30943> A_IWL<30942> A_IWL<30941> A_IWL<30940> A_IWL<30939> A_IWL<30938> A_IWL<30937> A_IWL<30936> A_IWL<30935> A_IWL<30934> A_IWL<30933> A_IWL<30932> A_IWL<30931> A_IWL<30930> A_IWL<30929> A_IWL<30928> A_IWL<30927> A_IWL<30926> A_IWL<30925> A_IWL<30924> A_IWL<30923> A_IWL<30922> A_IWL<30921> A_IWL<30920> A_IWL<30919> A_IWL<30918> A_IWL<30917> A_IWL<30916> A_IWL<30915> A_IWL<30914> A_IWL<30913> A_IWL<30912> A_IWL<30911> A_IWL<30910> A_IWL<30909> A_IWL<30908> A_IWL<30907> A_IWL<30906> A_IWL<30905> A_IWL<30904> A_IWL<30903> A_IWL<30902> A_IWL<30901> A_IWL<30900> A_IWL<30899> A_IWL<30898> A_IWL<30897> A_IWL<30896> A_IWL<30895> A_IWL<30894> A_IWL<30893> A_IWL<30892> A_IWL<30891> A_IWL<30890> A_IWL<30889> A_IWL<30888> A_IWL<30887> A_IWL<30886> A_IWL<30885> A_IWL<30884> A_IWL<30883> A_IWL<30882> A_IWL<30881> A_IWL<30880> A_IWL<30879> A_IWL<30878> A_IWL<30877> A_IWL<30876> A_IWL<30875> A_IWL<30874> A_IWL<30873> A_IWL<30872> A_IWL<30871> A_IWL<30870> A_IWL<30869> A_IWL<30868> A_IWL<30867> A_IWL<30866> A_IWL<30865> A_IWL<30864> A_IWL<30863> A_IWL<30862> A_IWL<30861> A_IWL<30860> A_IWL<30859> A_IWL<30858> A_IWL<30857> A_IWL<30856> A_IWL<30855> A_IWL<30854> A_IWL<30853> A_IWL<30852> A_IWL<30851> A_IWL<30850> A_IWL<30849> A_IWL<30848> A_IWL<30847> A_IWL<30846> A_IWL<30845> A_IWL<30844> A_IWL<30843> A_IWL<30842> A_IWL<30841> A_IWL<30840> A_IWL<30839> A_IWL<30838> A_IWL<30837> A_IWL<30836> A_IWL<30835> A_IWL<30834> A_IWL<30833> A_IWL<30832> A_IWL<30831> A_IWL<30830> A_IWL<30829> A_IWL<30828> A_IWL<30827> A_IWL<30826> A_IWL<30825> A_IWL<30824> A_IWL<30823> A_IWL<30822> A_IWL<30821> A_IWL<30820> A_IWL<30819> A_IWL<30818> A_IWL<30817> A_IWL<30816> A_IWL<30815> A_IWL<30814> A_IWL<30813> A_IWL<30812> A_IWL<30811> A_IWL<30810> A_IWL<30809> A_IWL<30808> A_IWL<30807> A_IWL<30806> A_IWL<30805> A_IWL<30804> A_IWL<30803> A_IWL<30802> A_IWL<30801> A_IWL<30800> A_IWL<30799> A_IWL<30798> A_IWL<30797> A_IWL<30796> A_IWL<30795> A_IWL<30794> A_IWL<30793> A_IWL<30792> A_IWL<30791> A_IWL<30790> A_IWL<30789> A_IWL<30788> A_IWL<30787> A_IWL<30786> A_IWL<30785> A_IWL<30784> A_IWL<30783> A_IWL<30782> A_IWL<30781> A_IWL<30780> A_IWL<30779> A_IWL<30778> A_IWL<30777> A_IWL<30776> A_IWL<30775> A_IWL<30774> A_IWL<30773> A_IWL<30772> A_IWL<30771> A_IWL<30770> A_IWL<30769> A_IWL<30768> A_IWL<30767> A_IWL<30766> A_IWL<30765> A_IWL<30764> A_IWL<30763> A_IWL<30762> A_IWL<30761> A_IWL<30760> A_IWL<30759> A_IWL<30758> A_IWL<30757> A_IWL<30756> A_IWL<30755> A_IWL<30754> A_IWL<30753> A_IWL<30752> A_IWL<30751> A_IWL<30750> A_IWL<30749> A_IWL<30748> A_IWL<30747> A_IWL<30746> A_IWL<30745> A_IWL<30744> A_IWL<30743> A_IWL<30742> A_IWL<30741> A_IWL<30740> A_IWL<30739> A_IWL<30738> A_IWL<30737> A_IWL<30736> A_IWL<30735> A_IWL<30734> A_IWL<30733> A_IWL<30732> A_IWL<30731> A_IWL<30730> A_IWL<30729> A_IWL<30728> A_IWL<30727> A_IWL<30726> A_IWL<30725> A_IWL<30724> A_IWL<30723> A_IWL<30722> A_IWL<30721> A_IWL<30720> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<59> A_BLC<119> A_BLC<118> A_BLC_TOP<119> A_BLC_TOP<118> A_BLT<119> A_BLT<118> A_BLT_TOP<119> A_BLT_TOP<118> A_IWL<30207> A_IWL<30206> A_IWL<30205> A_IWL<30204> A_IWL<30203> A_IWL<30202> A_IWL<30201> A_IWL<30200> A_IWL<30199> A_IWL<30198> A_IWL<30197> A_IWL<30196> A_IWL<30195> A_IWL<30194> A_IWL<30193> A_IWL<30192> A_IWL<30191> A_IWL<30190> A_IWL<30189> A_IWL<30188> A_IWL<30187> A_IWL<30186> A_IWL<30185> A_IWL<30184> A_IWL<30183> A_IWL<30182> A_IWL<30181> A_IWL<30180> A_IWL<30179> A_IWL<30178> A_IWL<30177> A_IWL<30176> A_IWL<30175> A_IWL<30174> A_IWL<30173> A_IWL<30172> A_IWL<30171> A_IWL<30170> A_IWL<30169> A_IWL<30168> A_IWL<30167> A_IWL<30166> A_IWL<30165> A_IWL<30164> A_IWL<30163> A_IWL<30162> A_IWL<30161> A_IWL<30160> A_IWL<30159> A_IWL<30158> A_IWL<30157> A_IWL<30156> A_IWL<30155> A_IWL<30154> A_IWL<30153> A_IWL<30152> A_IWL<30151> A_IWL<30150> A_IWL<30149> A_IWL<30148> A_IWL<30147> A_IWL<30146> A_IWL<30145> A_IWL<30144> A_IWL<30143> A_IWL<30142> A_IWL<30141> A_IWL<30140> A_IWL<30139> A_IWL<30138> A_IWL<30137> A_IWL<30136> A_IWL<30135> A_IWL<30134> A_IWL<30133> A_IWL<30132> A_IWL<30131> A_IWL<30130> A_IWL<30129> A_IWL<30128> A_IWL<30127> A_IWL<30126> A_IWL<30125> A_IWL<30124> A_IWL<30123> A_IWL<30122> A_IWL<30121> A_IWL<30120> A_IWL<30119> A_IWL<30118> A_IWL<30117> A_IWL<30116> A_IWL<30115> A_IWL<30114> A_IWL<30113> A_IWL<30112> A_IWL<30111> A_IWL<30110> A_IWL<30109> A_IWL<30108> A_IWL<30107> A_IWL<30106> A_IWL<30105> A_IWL<30104> A_IWL<30103> A_IWL<30102> A_IWL<30101> A_IWL<30100> A_IWL<30099> A_IWL<30098> A_IWL<30097> A_IWL<30096> A_IWL<30095> A_IWL<30094> A_IWL<30093> A_IWL<30092> A_IWL<30091> A_IWL<30090> A_IWL<30089> A_IWL<30088> A_IWL<30087> A_IWL<30086> A_IWL<30085> A_IWL<30084> A_IWL<30083> A_IWL<30082> A_IWL<30081> A_IWL<30080> A_IWL<30079> A_IWL<30078> A_IWL<30077> A_IWL<30076> A_IWL<30075> A_IWL<30074> A_IWL<30073> A_IWL<30072> A_IWL<30071> A_IWL<30070> A_IWL<30069> A_IWL<30068> A_IWL<30067> A_IWL<30066> A_IWL<30065> A_IWL<30064> A_IWL<30063> A_IWL<30062> A_IWL<30061> A_IWL<30060> A_IWL<30059> A_IWL<30058> A_IWL<30057> A_IWL<30056> A_IWL<30055> A_IWL<30054> A_IWL<30053> A_IWL<30052> A_IWL<30051> A_IWL<30050> A_IWL<30049> A_IWL<30048> A_IWL<30047> A_IWL<30046> A_IWL<30045> A_IWL<30044> A_IWL<30043> A_IWL<30042> A_IWL<30041> A_IWL<30040> A_IWL<30039> A_IWL<30038> A_IWL<30037> A_IWL<30036> A_IWL<30035> A_IWL<30034> A_IWL<30033> A_IWL<30032> A_IWL<30031> A_IWL<30030> A_IWL<30029> A_IWL<30028> A_IWL<30027> A_IWL<30026> A_IWL<30025> A_IWL<30024> A_IWL<30023> A_IWL<30022> A_IWL<30021> A_IWL<30020> A_IWL<30019> A_IWL<30018> A_IWL<30017> A_IWL<30016> A_IWL<30015> A_IWL<30014> A_IWL<30013> A_IWL<30012> A_IWL<30011> A_IWL<30010> A_IWL<30009> A_IWL<30008> A_IWL<30007> A_IWL<30006> A_IWL<30005> A_IWL<30004> A_IWL<30003> A_IWL<30002> A_IWL<30001> A_IWL<30000> A_IWL<29999> A_IWL<29998> A_IWL<29997> A_IWL<29996> A_IWL<29995> A_IWL<29994> A_IWL<29993> A_IWL<29992> A_IWL<29991> A_IWL<29990> A_IWL<29989> A_IWL<29988> A_IWL<29987> A_IWL<29986> A_IWL<29985> A_IWL<29984> A_IWL<29983> A_IWL<29982> A_IWL<29981> A_IWL<29980> A_IWL<29979> A_IWL<29978> A_IWL<29977> A_IWL<29976> A_IWL<29975> A_IWL<29974> A_IWL<29973> A_IWL<29972> A_IWL<29971> A_IWL<29970> A_IWL<29969> A_IWL<29968> A_IWL<29967> A_IWL<29966> A_IWL<29965> A_IWL<29964> A_IWL<29963> A_IWL<29962> A_IWL<29961> A_IWL<29960> A_IWL<29959> A_IWL<29958> A_IWL<29957> A_IWL<29956> A_IWL<29955> A_IWL<29954> A_IWL<29953> A_IWL<29952> A_IWL<29951> A_IWL<29950> A_IWL<29949> A_IWL<29948> A_IWL<29947> A_IWL<29946> A_IWL<29945> A_IWL<29944> A_IWL<29943> A_IWL<29942> A_IWL<29941> A_IWL<29940> A_IWL<29939> A_IWL<29938> A_IWL<29937> A_IWL<29936> A_IWL<29935> A_IWL<29934> A_IWL<29933> A_IWL<29932> A_IWL<29931> A_IWL<29930> A_IWL<29929> A_IWL<29928> A_IWL<29927> A_IWL<29926> A_IWL<29925> A_IWL<29924> A_IWL<29923> A_IWL<29922> A_IWL<29921> A_IWL<29920> A_IWL<29919> A_IWL<29918> A_IWL<29917> A_IWL<29916> A_IWL<29915> A_IWL<29914> A_IWL<29913> A_IWL<29912> A_IWL<29911> A_IWL<29910> A_IWL<29909> A_IWL<29908> A_IWL<29907> A_IWL<29906> A_IWL<29905> A_IWL<29904> A_IWL<29903> A_IWL<29902> A_IWL<29901> A_IWL<29900> A_IWL<29899> A_IWL<29898> A_IWL<29897> A_IWL<29896> A_IWL<29895> A_IWL<29894> A_IWL<29893> A_IWL<29892> A_IWL<29891> A_IWL<29890> A_IWL<29889> A_IWL<29888> A_IWL<29887> A_IWL<29886> A_IWL<29885> A_IWL<29884> A_IWL<29883> A_IWL<29882> A_IWL<29881> A_IWL<29880> A_IWL<29879> A_IWL<29878> A_IWL<29877> A_IWL<29876> A_IWL<29875> A_IWL<29874> A_IWL<29873> A_IWL<29872> A_IWL<29871> A_IWL<29870> A_IWL<29869> A_IWL<29868> A_IWL<29867> A_IWL<29866> A_IWL<29865> A_IWL<29864> A_IWL<29863> A_IWL<29862> A_IWL<29861> A_IWL<29860> A_IWL<29859> A_IWL<29858> A_IWL<29857> A_IWL<29856> A_IWL<29855> A_IWL<29854> A_IWL<29853> A_IWL<29852> A_IWL<29851> A_IWL<29850> A_IWL<29849> A_IWL<29848> A_IWL<29847> A_IWL<29846> A_IWL<29845> A_IWL<29844> A_IWL<29843> A_IWL<29842> A_IWL<29841> A_IWL<29840> A_IWL<29839> A_IWL<29838> A_IWL<29837> A_IWL<29836> A_IWL<29835> A_IWL<29834> A_IWL<29833> A_IWL<29832> A_IWL<29831> A_IWL<29830> A_IWL<29829> A_IWL<29828> A_IWL<29827> A_IWL<29826> A_IWL<29825> A_IWL<29824> A_IWL<29823> A_IWL<29822> A_IWL<29821> A_IWL<29820> A_IWL<29819> A_IWL<29818> A_IWL<29817> A_IWL<29816> A_IWL<29815> A_IWL<29814> A_IWL<29813> A_IWL<29812> A_IWL<29811> A_IWL<29810> A_IWL<29809> A_IWL<29808> A_IWL<29807> A_IWL<29806> A_IWL<29805> A_IWL<29804> A_IWL<29803> A_IWL<29802> A_IWL<29801> A_IWL<29800> A_IWL<29799> A_IWL<29798> A_IWL<29797> A_IWL<29796> A_IWL<29795> A_IWL<29794> A_IWL<29793> A_IWL<29792> A_IWL<29791> A_IWL<29790> A_IWL<29789> A_IWL<29788> A_IWL<29787> A_IWL<29786> A_IWL<29785> A_IWL<29784> A_IWL<29783> A_IWL<29782> A_IWL<29781> A_IWL<29780> A_IWL<29779> A_IWL<29778> A_IWL<29777> A_IWL<29776> A_IWL<29775> A_IWL<29774> A_IWL<29773> A_IWL<29772> A_IWL<29771> A_IWL<29770> A_IWL<29769> A_IWL<29768> A_IWL<29767> A_IWL<29766> A_IWL<29765> A_IWL<29764> A_IWL<29763> A_IWL<29762> A_IWL<29761> A_IWL<29760> A_IWL<29759> A_IWL<29758> A_IWL<29757> A_IWL<29756> A_IWL<29755> A_IWL<29754> A_IWL<29753> A_IWL<29752> A_IWL<29751> A_IWL<29750> A_IWL<29749> A_IWL<29748> A_IWL<29747> A_IWL<29746> A_IWL<29745> A_IWL<29744> A_IWL<29743> A_IWL<29742> A_IWL<29741> A_IWL<29740> A_IWL<29739> A_IWL<29738> A_IWL<29737> A_IWL<29736> A_IWL<29735> A_IWL<29734> A_IWL<29733> A_IWL<29732> A_IWL<29731> A_IWL<29730> A_IWL<29729> A_IWL<29728> A_IWL<29727> A_IWL<29726> A_IWL<29725> A_IWL<29724> A_IWL<29723> A_IWL<29722> A_IWL<29721> A_IWL<29720> A_IWL<29719> A_IWL<29718> A_IWL<29717> A_IWL<29716> A_IWL<29715> A_IWL<29714> A_IWL<29713> A_IWL<29712> A_IWL<29711> A_IWL<29710> A_IWL<29709> A_IWL<29708> A_IWL<29707> A_IWL<29706> A_IWL<29705> A_IWL<29704> A_IWL<29703> A_IWL<29702> A_IWL<29701> A_IWL<29700> A_IWL<29699> A_IWL<29698> A_IWL<29697> A_IWL<29696> A_IWL<30719> A_IWL<30718> A_IWL<30717> A_IWL<30716> A_IWL<30715> A_IWL<30714> A_IWL<30713> A_IWL<30712> A_IWL<30711> A_IWL<30710> A_IWL<30709> A_IWL<30708> A_IWL<30707> A_IWL<30706> A_IWL<30705> A_IWL<30704> A_IWL<30703> A_IWL<30702> A_IWL<30701> A_IWL<30700> A_IWL<30699> A_IWL<30698> A_IWL<30697> A_IWL<30696> A_IWL<30695> A_IWL<30694> A_IWL<30693> A_IWL<30692> A_IWL<30691> A_IWL<30690> A_IWL<30689> A_IWL<30688> A_IWL<30687> A_IWL<30686> A_IWL<30685> A_IWL<30684> A_IWL<30683> A_IWL<30682> A_IWL<30681> A_IWL<30680> A_IWL<30679> A_IWL<30678> A_IWL<30677> A_IWL<30676> A_IWL<30675> A_IWL<30674> A_IWL<30673> A_IWL<30672> A_IWL<30671> A_IWL<30670> A_IWL<30669> A_IWL<30668> A_IWL<30667> A_IWL<30666> A_IWL<30665> A_IWL<30664> A_IWL<30663> A_IWL<30662> A_IWL<30661> A_IWL<30660> A_IWL<30659> A_IWL<30658> A_IWL<30657> A_IWL<30656> A_IWL<30655> A_IWL<30654> A_IWL<30653> A_IWL<30652> A_IWL<30651> A_IWL<30650> A_IWL<30649> A_IWL<30648> A_IWL<30647> A_IWL<30646> A_IWL<30645> A_IWL<30644> A_IWL<30643> A_IWL<30642> A_IWL<30641> A_IWL<30640> A_IWL<30639> A_IWL<30638> A_IWL<30637> A_IWL<30636> A_IWL<30635> A_IWL<30634> A_IWL<30633> A_IWL<30632> A_IWL<30631> A_IWL<30630> A_IWL<30629> A_IWL<30628> A_IWL<30627> A_IWL<30626> A_IWL<30625> A_IWL<30624> A_IWL<30623> A_IWL<30622> A_IWL<30621> A_IWL<30620> A_IWL<30619> A_IWL<30618> A_IWL<30617> A_IWL<30616> A_IWL<30615> A_IWL<30614> A_IWL<30613> A_IWL<30612> A_IWL<30611> A_IWL<30610> A_IWL<30609> A_IWL<30608> A_IWL<30607> A_IWL<30606> A_IWL<30605> A_IWL<30604> A_IWL<30603> A_IWL<30602> A_IWL<30601> A_IWL<30600> A_IWL<30599> A_IWL<30598> A_IWL<30597> A_IWL<30596> A_IWL<30595> A_IWL<30594> A_IWL<30593> A_IWL<30592> A_IWL<30591> A_IWL<30590> A_IWL<30589> A_IWL<30588> A_IWL<30587> A_IWL<30586> A_IWL<30585> A_IWL<30584> A_IWL<30583> A_IWL<30582> A_IWL<30581> A_IWL<30580> A_IWL<30579> A_IWL<30578> A_IWL<30577> A_IWL<30576> A_IWL<30575> A_IWL<30574> A_IWL<30573> A_IWL<30572> A_IWL<30571> A_IWL<30570> A_IWL<30569> A_IWL<30568> A_IWL<30567> A_IWL<30566> A_IWL<30565> A_IWL<30564> A_IWL<30563> A_IWL<30562> A_IWL<30561> A_IWL<30560> A_IWL<30559> A_IWL<30558> A_IWL<30557> A_IWL<30556> A_IWL<30555> A_IWL<30554> A_IWL<30553> A_IWL<30552> A_IWL<30551> A_IWL<30550> A_IWL<30549> A_IWL<30548> A_IWL<30547> A_IWL<30546> A_IWL<30545> A_IWL<30544> A_IWL<30543> A_IWL<30542> A_IWL<30541> A_IWL<30540> A_IWL<30539> A_IWL<30538> A_IWL<30537> A_IWL<30536> A_IWL<30535> A_IWL<30534> A_IWL<30533> A_IWL<30532> A_IWL<30531> A_IWL<30530> A_IWL<30529> A_IWL<30528> A_IWL<30527> A_IWL<30526> A_IWL<30525> A_IWL<30524> A_IWL<30523> A_IWL<30522> A_IWL<30521> A_IWL<30520> A_IWL<30519> A_IWL<30518> A_IWL<30517> A_IWL<30516> A_IWL<30515> A_IWL<30514> A_IWL<30513> A_IWL<30512> A_IWL<30511> A_IWL<30510> A_IWL<30509> A_IWL<30508> A_IWL<30507> A_IWL<30506> A_IWL<30505> A_IWL<30504> A_IWL<30503> A_IWL<30502> A_IWL<30501> A_IWL<30500> A_IWL<30499> A_IWL<30498> A_IWL<30497> A_IWL<30496> A_IWL<30495> A_IWL<30494> A_IWL<30493> A_IWL<30492> A_IWL<30491> A_IWL<30490> A_IWL<30489> A_IWL<30488> A_IWL<30487> A_IWL<30486> A_IWL<30485> A_IWL<30484> A_IWL<30483> A_IWL<30482> A_IWL<30481> A_IWL<30480> A_IWL<30479> A_IWL<30478> A_IWL<30477> A_IWL<30476> A_IWL<30475> A_IWL<30474> A_IWL<30473> A_IWL<30472> A_IWL<30471> A_IWL<30470> A_IWL<30469> A_IWL<30468> A_IWL<30467> A_IWL<30466> A_IWL<30465> A_IWL<30464> A_IWL<30463> A_IWL<30462> A_IWL<30461> A_IWL<30460> A_IWL<30459> A_IWL<30458> A_IWL<30457> A_IWL<30456> A_IWL<30455> A_IWL<30454> A_IWL<30453> A_IWL<30452> A_IWL<30451> A_IWL<30450> A_IWL<30449> A_IWL<30448> A_IWL<30447> A_IWL<30446> A_IWL<30445> A_IWL<30444> A_IWL<30443> A_IWL<30442> A_IWL<30441> A_IWL<30440> A_IWL<30439> A_IWL<30438> A_IWL<30437> A_IWL<30436> A_IWL<30435> A_IWL<30434> A_IWL<30433> A_IWL<30432> A_IWL<30431> A_IWL<30430> A_IWL<30429> A_IWL<30428> A_IWL<30427> A_IWL<30426> A_IWL<30425> A_IWL<30424> A_IWL<30423> A_IWL<30422> A_IWL<30421> A_IWL<30420> A_IWL<30419> A_IWL<30418> A_IWL<30417> A_IWL<30416> A_IWL<30415> A_IWL<30414> A_IWL<30413> A_IWL<30412> A_IWL<30411> A_IWL<30410> A_IWL<30409> A_IWL<30408> A_IWL<30407> A_IWL<30406> A_IWL<30405> A_IWL<30404> A_IWL<30403> A_IWL<30402> A_IWL<30401> A_IWL<30400> A_IWL<30399> A_IWL<30398> A_IWL<30397> A_IWL<30396> A_IWL<30395> A_IWL<30394> A_IWL<30393> A_IWL<30392> A_IWL<30391> A_IWL<30390> A_IWL<30389> A_IWL<30388> A_IWL<30387> A_IWL<30386> A_IWL<30385> A_IWL<30384> A_IWL<30383> A_IWL<30382> A_IWL<30381> A_IWL<30380> A_IWL<30379> A_IWL<30378> A_IWL<30377> A_IWL<30376> A_IWL<30375> A_IWL<30374> A_IWL<30373> A_IWL<30372> A_IWL<30371> A_IWL<30370> A_IWL<30369> A_IWL<30368> A_IWL<30367> A_IWL<30366> A_IWL<30365> A_IWL<30364> A_IWL<30363> A_IWL<30362> A_IWL<30361> A_IWL<30360> A_IWL<30359> A_IWL<30358> A_IWL<30357> A_IWL<30356> A_IWL<30355> A_IWL<30354> A_IWL<30353> A_IWL<30352> A_IWL<30351> A_IWL<30350> A_IWL<30349> A_IWL<30348> A_IWL<30347> A_IWL<30346> A_IWL<30345> A_IWL<30344> A_IWL<30343> A_IWL<30342> A_IWL<30341> A_IWL<30340> A_IWL<30339> A_IWL<30338> A_IWL<30337> A_IWL<30336> A_IWL<30335> A_IWL<30334> A_IWL<30333> A_IWL<30332> A_IWL<30331> A_IWL<30330> A_IWL<30329> A_IWL<30328> A_IWL<30327> A_IWL<30326> A_IWL<30325> A_IWL<30324> A_IWL<30323> A_IWL<30322> A_IWL<30321> A_IWL<30320> A_IWL<30319> A_IWL<30318> A_IWL<30317> A_IWL<30316> A_IWL<30315> A_IWL<30314> A_IWL<30313> A_IWL<30312> A_IWL<30311> A_IWL<30310> A_IWL<30309> A_IWL<30308> A_IWL<30307> A_IWL<30306> A_IWL<30305> A_IWL<30304> A_IWL<30303> A_IWL<30302> A_IWL<30301> A_IWL<30300> A_IWL<30299> A_IWL<30298> A_IWL<30297> A_IWL<30296> A_IWL<30295> A_IWL<30294> A_IWL<30293> A_IWL<30292> A_IWL<30291> A_IWL<30290> A_IWL<30289> A_IWL<30288> A_IWL<30287> A_IWL<30286> A_IWL<30285> A_IWL<30284> A_IWL<30283> A_IWL<30282> A_IWL<30281> A_IWL<30280> A_IWL<30279> A_IWL<30278> A_IWL<30277> A_IWL<30276> A_IWL<30275> A_IWL<30274> A_IWL<30273> A_IWL<30272> A_IWL<30271> A_IWL<30270> A_IWL<30269> A_IWL<30268> A_IWL<30267> A_IWL<30266> A_IWL<30265> A_IWL<30264> A_IWL<30263> A_IWL<30262> A_IWL<30261> A_IWL<30260> A_IWL<30259> A_IWL<30258> A_IWL<30257> A_IWL<30256> A_IWL<30255> A_IWL<30254> A_IWL<30253> A_IWL<30252> A_IWL<30251> A_IWL<30250> A_IWL<30249> A_IWL<30248> A_IWL<30247> A_IWL<30246> A_IWL<30245> A_IWL<30244> A_IWL<30243> A_IWL<30242> A_IWL<30241> A_IWL<30240> A_IWL<30239> A_IWL<30238> A_IWL<30237> A_IWL<30236> A_IWL<30235> A_IWL<30234> A_IWL<30233> A_IWL<30232> A_IWL<30231> A_IWL<30230> A_IWL<30229> A_IWL<30228> A_IWL<30227> A_IWL<30226> A_IWL<30225> A_IWL<30224> A_IWL<30223> A_IWL<30222> A_IWL<30221> A_IWL<30220> A_IWL<30219> A_IWL<30218> A_IWL<30217> A_IWL<30216> A_IWL<30215> A_IWL<30214> A_IWL<30213> A_IWL<30212> A_IWL<30211> A_IWL<30210> A_IWL<30209> A_IWL<30208> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<58> A_BLC<117> A_BLC<116> A_BLC_TOP<117> A_BLC_TOP<116> A_BLT<117> A_BLT<116> A_BLT_TOP<117> A_BLT_TOP<116> A_IWL<29695> A_IWL<29694> A_IWL<29693> A_IWL<29692> A_IWL<29691> A_IWL<29690> A_IWL<29689> A_IWL<29688> A_IWL<29687> A_IWL<29686> A_IWL<29685> A_IWL<29684> A_IWL<29683> A_IWL<29682> A_IWL<29681> A_IWL<29680> A_IWL<29679> A_IWL<29678> A_IWL<29677> A_IWL<29676> A_IWL<29675> A_IWL<29674> A_IWL<29673> A_IWL<29672> A_IWL<29671> A_IWL<29670> A_IWL<29669> A_IWL<29668> A_IWL<29667> A_IWL<29666> A_IWL<29665> A_IWL<29664> A_IWL<29663> A_IWL<29662> A_IWL<29661> A_IWL<29660> A_IWL<29659> A_IWL<29658> A_IWL<29657> A_IWL<29656> A_IWL<29655> A_IWL<29654> A_IWL<29653> A_IWL<29652> A_IWL<29651> A_IWL<29650> A_IWL<29649> A_IWL<29648> A_IWL<29647> A_IWL<29646> A_IWL<29645> A_IWL<29644> A_IWL<29643> A_IWL<29642> A_IWL<29641> A_IWL<29640> A_IWL<29639> A_IWL<29638> A_IWL<29637> A_IWL<29636> A_IWL<29635> A_IWL<29634> A_IWL<29633> A_IWL<29632> A_IWL<29631> A_IWL<29630> A_IWL<29629> A_IWL<29628> A_IWL<29627> A_IWL<29626> A_IWL<29625> A_IWL<29624> A_IWL<29623> A_IWL<29622> A_IWL<29621> A_IWL<29620> A_IWL<29619> A_IWL<29618> A_IWL<29617> A_IWL<29616> A_IWL<29615> A_IWL<29614> A_IWL<29613> A_IWL<29612> A_IWL<29611> A_IWL<29610> A_IWL<29609> A_IWL<29608> A_IWL<29607> A_IWL<29606> A_IWL<29605> A_IWL<29604> A_IWL<29603> A_IWL<29602> A_IWL<29601> A_IWL<29600> A_IWL<29599> A_IWL<29598> A_IWL<29597> A_IWL<29596> A_IWL<29595> A_IWL<29594> A_IWL<29593> A_IWL<29592> A_IWL<29591> A_IWL<29590> A_IWL<29589> A_IWL<29588> A_IWL<29587> A_IWL<29586> A_IWL<29585> A_IWL<29584> A_IWL<29583> A_IWL<29582> A_IWL<29581> A_IWL<29580> A_IWL<29579> A_IWL<29578> A_IWL<29577> A_IWL<29576> A_IWL<29575> A_IWL<29574> A_IWL<29573> A_IWL<29572> A_IWL<29571> A_IWL<29570> A_IWL<29569> A_IWL<29568> A_IWL<29567> A_IWL<29566> A_IWL<29565> A_IWL<29564> A_IWL<29563> A_IWL<29562> A_IWL<29561> A_IWL<29560> A_IWL<29559> A_IWL<29558> A_IWL<29557> A_IWL<29556> A_IWL<29555> A_IWL<29554> A_IWL<29553> A_IWL<29552> A_IWL<29551> A_IWL<29550> A_IWL<29549> A_IWL<29548> A_IWL<29547> A_IWL<29546> A_IWL<29545> A_IWL<29544> A_IWL<29543> A_IWL<29542> A_IWL<29541> A_IWL<29540> A_IWL<29539> A_IWL<29538> A_IWL<29537> A_IWL<29536> A_IWL<29535> A_IWL<29534> A_IWL<29533> A_IWL<29532> A_IWL<29531> A_IWL<29530> A_IWL<29529> A_IWL<29528> A_IWL<29527> A_IWL<29526> A_IWL<29525> A_IWL<29524> A_IWL<29523> A_IWL<29522> A_IWL<29521> A_IWL<29520> A_IWL<29519> A_IWL<29518> A_IWL<29517> A_IWL<29516> A_IWL<29515> A_IWL<29514> A_IWL<29513> A_IWL<29512> A_IWL<29511> A_IWL<29510> A_IWL<29509> A_IWL<29508> A_IWL<29507> A_IWL<29506> A_IWL<29505> A_IWL<29504> A_IWL<29503> A_IWL<29502> A_IWL<29501> A_IWL<29500> A_IWL<29499> A_IWL<29498> A_IWL<29497> A_IWL<29496> A_IWL<29495> A_IWL<29494> A_IWL<29493> A_IWL<29492> A_IWL<29491> A_IWL<29490> A_IWL<29489> A_IWL<29488> A_IWL<29487> A_IWL<29486> A_IWL<29485> A_IWL<29484> A_IWL<29483> A_IWL<29482> A_IWL<29481> A_IWL<29480> A_IWL<29479> A_IWL<29478> A_IWL<29477> A_IWL<29476> A_IWL<29475> A_IWL<29474> A_IWL<29473> A_IWL<29472> A_IWL<29471> A_IWL<29470> A_IWL<29469> A_IWL<29468> A_IWL<29467> A_IWL<29466> A_IWL<29465> A_IWL<29464> A_IWL<29463> A_IWL<29462> A_IWL<29461> A_IWL<29460> A_IWL<29459> A_IWL<29458> A_IWL<29457> A_IWL<29456> A_IWL<29455> A_IWL<29454> A_IWL<29453> A_IWL<29452> A_IWL<29451> A_IWL<29450> A_IWL<29449> A_IWL<29448> A_IWL<29447> A_IWL<29446> A_IWL<29445> A_IWL<29444> A_IWL<29443> A_IWL<29442> A_IWL<29441> A_IWL<29440> A_IWL<29439> A_IWL<29438> A_IWL<29437> A_IWL<29436> A_IWL<29435> A_IWL<29434> A_IWL<29433> A_IWL<29432> A_IWL<29431> A_IWL<29430> A_IWL<29429> A_IWL<29428> A_IWL<29427> A_IWL<29426> A_IWL<29425> A_IWL<29424> A_IWL<29423> A_IWL<29422> A_IWL<29421> A_IWL<29420> A_IWL<29419> A_IWL<29418> A_IWL<29417> A_IWL<29416> A_IWL<29415> A_IWL<29414> A_IWL<29413> A_IWL<29412> A_IWL<29411> A_IWL<29410> A_IWL<29409> A_IWL<29408> A_IWL<29407> A_IWL<29406> A_IWL<29405> A_IWL<29404> A_IWL<29403> A_IWL<29402> A_IWL<29401> A_IWL<29400> A_IWL<29399> A_IWL<29398> A_IWL<29397> A_IWL<29396> A_IWL<29395> A_IWL<29394> A_IWL<29393> A_IWL<29392> A_IWL<29391> A_IWL<29390> A_IWL<29389> A_IWL<29388> A_IWL<29387> A_IWL<29386> A_IWL<29385> A_IWL<29384> A_IWL<29383> A_IWL<29382> A_IWL<29381> A_IWL<29380> A_IWL<29379> A_IWL<29378> A_IWL<29377> A_IWL<29376> A_IWL<29375> A_IWL<29374> A_IWL<29373> A_IWL<29372> A_IWL<29371> A_IWL<29370> A_IWL<29369> A_IWL<29368> A_IWL<29367> A_IWL<29366> A_IWL<29365> A_IWL<29364> A_IWL<29363> A_IWL<29362> A_IWL<29361> A_IWL<29360> A_IWL<29359> A_IWL<29358> A_IWL<29357> A_IWL<29356> A_IWL<29355> A_IWL<29354> A_IWL<29353> A_IWL<29352> A_IWL<29351> A_IWL<29350> A_IWL<29349> A_IWL<29348> A_IWL<29347> A_IWL<29346> A_IWL<29345> A_IWL<29344> A_IWL<29343> A_IWL<29342> A_IWL<29341> A_IWL<29340> A_IWL<29339> A_IWL<29338> A_IWL<29337> A_IWL<29336> A_IWL<29335> A_IWL<29334> A_IWL<29333> A_IWL<29332> A_IWL<29331> A_IWL<29330> A_IWL<29329> A_IWL<29328> A_IWL<29327> A_IWL<29326> A_IWL<29325> A_IWL<29324> A_IWL<29323> A_IWL<29322> A_IWL<29321> A_IWL<29320> A_IWL<29319> A_IWL<29318> A_IWL<29317> A_IWL<29316> A_IWL<29315> A_IWL<29314> A_IWL<29313> A_IWL<29312> A_IWL<29311> A_IWL<29310> A_IWL<29309> A_IWL<29308> A_IWL<29307> A_IWL<29306> A_IWL<29305> A_IWL<29304> A_IWL<29303> A_IWL<29302> A_IWL<29301> A_IWL<29300> A_IWL<29299> A_IWL<29298> A_IWL<29297> A_IWL<29296> A_IWL<29295> A_IWL<29294> A_IWL<29293> A_IWL<29292> A_IWL<29291> A_IWL<29290> A_IWL<29289> A_IWL<29288> A_IWL<29287> A_IWL<29286> A_IWL<29285> A_IWL<29284> A_IWL<29283> A_IWL<29282> A_IWL<29281> A_IWL<29280> A_IWL<29279> A_IWL<29278> A_IWL<29277> A_IWL<29276> A_IWL<29275> A_IWL<29274> A_IWL<29273> A_IWL<29272> A_IWL<29271> A_IWL<29270> A_IWL<29269> A_IWL<29268> A_IWL<29267> A_IWL<29266> A_IWL<29265> A_IWL<29264> A_IWL<29263> A_IWL<29262> A_IWL<29261> A_IWL<29260> A_IWL<29259> A_IWL<29258> A_IWL<29257> A_IWL<29256> A_IWL<29255> A_IWL<29254> A_IWL<29253> A_IWL<29252> A_IWL<29251> A_IWL<29250> A_IWL<29249> A_IWL<29248> A_IWL<29247> A_IWL<29246> A_IWL<29245> A_IWL<29244> A_IWL<29243> A_IWL<29242> A_IWL<29241> A_IWL<29240> A_IWL<29239> A_IWL<29238> A_IWL<29237> A_IWL<29236> A_IWL<29235> A_IWL<29234> A_IWL<29233> A_IWL<29232> A_IWL<29231> A_IWL<29230> A_IWL<29229> A_IWL<29228> A_IWL<29227> A_IWL<29226> A_IWL<29225> A_IWL<29224> A_IWL<29223> A_IWL<29222> A_IWL<29221> A_IWL<29220> A_IWL<29219> A_IWL<29218> A_IWL<29217> A_IWL<29216> A_IWL<29215> A_IWL<29214> A_IWL<29213> A_IWL<29212> A_IWL<29211> A_IWL<29210> A_IWL<29209> A_IWL<29208> A_IWL<29207> A_IWL<29206> A_IWL<29205> A_IWL<29204> A_IWL<29203> A_IWL<29202> A_IWL<29201> A_IWL<29200> A_IWL<29199> A_IWL<29198> A_IWL<29197> A_IWL<29196> A_IWL<29195> A_IWL<29194> A_IWL<29193> A_IWL<29192> A_IWL<29191> A_IWL<29190> A_IWL<29189> A_IWL<29188> A_IWL<29187> A_IWL<29186> A_IWL<29185> A_IWL<29184> A_IWL<30207> A_IWL<30206> A_IWL<30205> A_IWL<30204> A_IWL<30203> A_IWL<30202> A_IWL<30201> A_IWL<30200> A_IWL<30199> A_IWL<30198> A_IWL<30197> A_IWL<30196> A_IWL<30195> A_IWL<30194> A_IWL<30193> A_IWL<30192> A_IWL<30191> A_IWL<30190> A_IWL<30189> A_IWL<30188> A_IWL<30187> A_IWL<30186> A_IWL<30185> A_IWL<30184> A_IWL<30183> A_IWL<30182> A_IWL<30181> A_IWL<30180> A_IWL<30179> A_IWL<30178> A_IWL<30177> A_IWL<30176> A_IWL<30175> A_IWL<30174> A_IWL<30173> A_IWL<30172> A_IWL<30171> A_IWL<30170> A_IWL<30169> A_IWL<30168> A_IWL<30167> A_IWL<30166> A_IWL<30165> A_IWL<30164> A_IWL<30163> A_IWL<30162> A_IWL<30161> A_IWL<30160> A_IWL<30159> A_IWL<30158> A_IWL<30157> A_IWL<30156> A_IWL<30155> A_IWL<30154> A_IWL<30153> A_IWL<30152> A_IWL<30151> A_IWL<30150> A_IWL<30149> A_IWL<30148> A_IWL<30147> A_IWL<30146> A_IWL<30145> A_IWL<30144> A_IWL<30143> A_IWL<30142> A_IWL<30141> A_IWL<30140> A_IWL<30139> A_IWL<30138> A_IWL<30137> A_IWL<30136> A_IWL<30135> A_IWL<30134> A_IWL<30133> A_IWL<30132> A_IWL<30131> A_IWL<30130> A_IWL<30129> A_IWL<30128> A_IWL<30127> A_IWL<30126> A_IWL<30125> A_IWL<30124> A_IWL<30123> A_IWL<30122> A_IWL<30121> A_IWL<30120> A_IWL<30119> A_IWL<30118> A_IWL<30117> A_IWL<30116> A_IWL<30115> A_IWL<30114> A_IWL<30113> A_IWL<30112> A_IWL<30111> A_IWL<30110> A_IWL<30109> A_IWL<30108> A_IWL<30107> A_IWL<30106> A_IWL<30105> A_IWL<30104> A_IWL<30103> A_IWL<30102> A_IWL<30101> A_IWL<30100> A_IWL<30099> A_IWL<30098> A_IWL<30097> A_IWL<30096> A_IWL<30095> A_IWL<30094> A_IWL<30093> A_IWL<30092> A_IWL<30091> A_IWL<30090> A_IWL<30089> A_IWL<30088> A_IWL<30087> A_IWL<30086> A_IWL<30085> A_IWL<30084> A_IWL<30083> A_IWL<30082> A_IWL<30081> A_IWL<30080> A_IWL<30079> A_IWL<30078> A_IWL<30077> A_IWL<30076> A_IWL<30075> A_IWL<30074> A_IWL<30073> A_IWL<30072> A_IWL<30071> A_IWL<30070> A_IWL<30069> A_IWL<30068> A_IWL<30067> A_IWL<30066> A_IWL<30065> A_IWL<30064> A_IWL<30063> A_IWL<30062> A_IWL<30061> A_IWL<30060> A_IWL<30059> A_IWL<30058> A_IWL<30057> A_IWL<30056> A_IWL<30055> A_IWL<30054> A_IWL<30053> A_IWL<30052> A_IWL<30051> A_IWL<30050> A_IWL<30049> A_IWL<30048> A_IWL<30047> A_IWL<30046> A_IWL<30045> A_IWL<30044> A_IWL<30043> A_IWL<30042> A_IWL<30041> A_IWL<30040> A_IWL<30039> A_IWL<30038> A_IWL<30037> A_IWL<30036> A_IWL<30035> A_IWL<30034> A_IWL<30033> A_IWL<30032> A_IWL<30031> A_IWL<30030> A_IWL<30029> A_IWL<30028> A_IWL<30027> A_IWL<30026> A_IWL<30025> A_IWL<30024> A_IWL<30023> A_IWL<30022> A_IWL<30021> A_IWL<30020> A_IWL<30019> A_IWL<30018> A_IWL<30017> A_IWL<30016> A_IWL<30015> A_IWL<30014> A_IWL<30013> A_IWL<30012> A_IWL<30011> A_IWL<30010> A_IWL<30009> A_IWL<30008> A_IWL<30007> A_IWL<30006> A_IWL<30005> A_IWL<30004> A_IWL<30003> A_IWL<30002> A_IWL<30001> A_IWL<30000> A_IWL<29999> A_IWL<29998> A_IWL<29997> A_IWL<29996> A_IWL<29995> A_IWL<29994> A_IWL<29993> A_IWL<29992> A_IWL<29991> A_IWL<29990> A_IWL<29989> A_IWL<29988> A_IWL<29987> A_IWL<29986> A_IWL<29985> A_IWL<29984> A_IWL<29983> A_IWL<29982> A_IWL<29981> A_IWL<29980> A_IWL<29979> A_IWL<29978> A_IWL<29977> A_IWL<29976> A_IWL<29975> A_IWL<29974> A_IWL<29973> A_IWL<29972> A_IWL<29971> A_IWL<29970> A_IWL<29969> A_IWL<29968> A_IWL<29967> A_IWL<29966> A_IWL<29965> A_IWL<29964> A_IWL<29963> A_IWL<29962> A_IWL<29961> A_IWL<29960> A_IWL<29959> A_IWL<29958> A_IWL<29957> A_IWL<29956> A_IWL<29955> A_IWL<29954> A_IWL<29953> A_IWL<29952> A_IWL<29951> A_IWL<29950> A_IWL<29949> A_IWL<29948> A_IWL<29947> A_IWL<29946> A_IWL<29945> A_IWL<29944> A_IWL<29943> A_IWL<29942> A_IWL<29941> A_IWL<29940> A_IWL<29939> A_IWL<29938> A_IWL<29937> A_IWL<29936> A_IWL<29935> A_IWL<29934> A_IWL<29933> A_IWL<29932> A_IWL<29931> A_IWL<29930> A_IWL<29929> A_IWL<29928> A_IWL<29927> A_IWL<29926> A_IWL<29925> A_IWL<29924> A_IWL<29923> A_IWL<29922> A_IWL<29921> A_IWL<29920> A_IWL<29919> A_IWL<29918> A_IWL<29917> A_IWL<29916> A_IWL<29915> A_IWL<29914> A_IWL<29913> A_IWL<29912> A_IWL<29911> A_IWL<29910> A_IWL<29909> A_IWL<29908> A_IWL<29907> A_IWL<29906> A_IWL<29905> A_IWL<29904> A_IWL<29903> A_IWL<29902> A_IWL<29901> A_IWL<29900> A_IWL<29899> A_IWL<29898> A_IWL<29897> A_IWL<29896> A_IWL<29895> A_IWL<29894> A_IWL<29893> A_IWL<29892> A_IWL<29891> A_IWL<29890> A_IWL<29889> A_IWL<29888> A_IWL<29887> A_IWL<29886> A_IWL<29885> A_IWL<29884> A_IWL<29883> A_IWL<29882> A_IWL<29881> A_IWL<29880> A_IWL<29879> A_IWL<29878> A_IWL<29877> A_IWL<29876> A_IWL<29875> A_IWL<29874> A_IWL<29873> A_IWL<29872> A_IWL<29871> A_IWL<29870> A_IWL<29869> A_IWL<29868> A_IWL<29867> A_IWL<29866> A_IWL<29865> A_IWL<29864> A_IWL<29863> A_IWL<29862> A_IWL<29861> A_IWL<29860> A_IWL<29859> A_IWL<29858> A_IWL<29857> A_IWL<29856> A_IWL<29855> A_IWL<29854> A_IWL<29853> A_IWL<29852> A_IWL<29851> A_IWL<29850> A_IWL<29849> A_IWL<29848> A_IWL<29847> A_IWL<29846> A_IWL<29845> A_IWL<29844> A_IWL<29843> A_IWL<29842> A_IWL<29841> A_IWL<29840> A_IWL<29839> A_IWL<29838> A_IWL<29837> A_IWL<29836> A_IWL<29835> A_IWL<29834> A_IWL<29833> A_IWL<29832> A_IWL<29831> A_IWL<29830> A_IWL<29829> A_IWL<29828> A_IWL<29827> A_IWL<29826> A_IWL<29825> A_IWL<29824> A_IWL<29823> A_IWL<29822> A_IWL<29821> A_IWL<29820> A_IWL<29819> A_IWL<29818> A_IWL<29817> A_IWL<29816> A_IWL<29815> A_IWL<29814> A_IWL<29813> A_IWL<29812> A_IWL<29811> A_IWL<29810> A_IWL<29809> A_IWL<29808> A_IWL<29807> A_IWL<29806> A_IWL<29805> A_IWL<29804> A_IWL<29803> A_IWL<29802> A_IWL<29801> A_IWL<29800> A_IWL<29799> A_IWL<29798> A_IWL<29797> A_IWL<29796> A_IWL<29795> A_IWL<29794> A_IWL<29793> A_IWL<29792> A_IWL<29791> A_IWL<29790> A_IWL<29789> A_IWL<29788> A_IWL<29787> A_IWL<29786> A_IWL<29785> A_IWL<29784> A_IWL<29783> A_IWL<29782> A_IWL<29781> A_IWL<29780> A_IWL<29779> A_IWL<29778> A_IWL<29777> A_IWL<29776> A_IWL<29775> A_IWL<29774> A_IWL<29773> A_IWL<29772> A_IWL<29771> A_IWL<29770> A_IWL<29769> A_IWL<29768> A_IWL<29767> A_IWL<29766> A_IWL<29765> A_IWL<29764> A_IWL<29763> A_IWL<29762> A_IWL<29761> A_IWL<29760> A_IWL<29759> A_IWL<29758> A_IWL<29757> A_IWL<29756> A_IWL<29755> A_IWL<29754> A_IWL<29753> A_IWL<29752> A_IWL<29751> A_IWL<29750> A_IWL<29749> A_IWL<29748> A_IWL<29747> A_IWL<29746> A_IWL<29745> A_IWL<29744> A_IWL<29743> A_IWL<29742> A_IWL<29741> A_IWL<29740> A_IWL<29739> A_IWL<29738> A_IWL<29737> A_IWL<29736> A_IWL<29735> A_IWL<29734> A_IWL<29733> A_IWL<29732> A_IWL<29731> A_IWL<29730> A_IWL<29729> A_IWL<29728> A_IWL<29727> A_IWL<29726> A_IWL<29725> A_IWL<29724> A_IWL<29723> A_IWL<29722> A_IWL<29721> A_IWL<29720> A_IWL<29719> A_IWL<29718> A_IWL<29717> A_IWL<29716> A_IWL<29715> A_IWL<29714> A_IWL<29713> A_IWL<29712> A_IWL<29711> A_IWL<29710> A_IWL<29709> A_IWL<29708> A_IWL<29707> A_IWL<29706> A_IWL<29705> A_IWL<29704> A_IWL<29703> A_IWL<29702> A_IWL<29701> A_IWL<29700> A_IWL<29699> A_IWL<29698> A_IWL<29697> A_IWL<29696> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<57> A_BLC<115> A_BLC<114> A_BLC_TOP<115> A_BLC_TOP<114> A_BLT<115> A_BLT<114> A_BLT_TOP<115> A_BLT_TOP<114> A_IWL<29183> A_IWL<29182> A_IWL<29181> A_IWL<29180> A_IWL<29179> A_IWL<29178> A_IWL<29177> A_IWL<29176> A_IWL<29175> A_IWL<29174> A_IWL<29173> A_IWL<29172> A_IWL<29171> A_IWL<29170> A_IWL<29169> A_IWL<29168> A_IWL<29167> A_IWL<29166> A_IWL<29165> A_IWL<29164> A_IWL<29163> A_IWL<29162> A_IWL<29161> A_IWL<29160> A_IWL<29159> A_IWL<29158> A_IWL<29157> A_IWL<29156> A_IWL<29155> A_IWL<29154> A_IWL<29153> A_IWL<29152> A_IWL<29151> A_IWL<29150> A_IWL<29149> A_IWL<29148> A_IWL<29147> A_IWL<29146> A_IWL<29145> A_IWL<29144> A_IWL<29143> A_IWL<29142> A_IWL<29141> A_IWL<29140> A_IWL<29139> A_IWL<29138> A_IWL<29137> A_IWL<29136> A_IWL<29135> A_IWL<29134> A_IWL<29133> A_IWL<29132> A_IWL<29131> A_IWL<29130> A_IWL<29129> A_IWL<29128> A_IWL<29127> A_IWL<29126> A_IWL<29125> A_IWL<29124> A_IWL<29123> A_IWL<29122> A_IWL<29121> A_IWL<29120> A_IWL<29119> A_IWL<29118> A_IWL<29117> A_IWL<29116> A_IWL<29115> A_IWL<29114> A_IWL<29113> A_IWL<29112> A_IWL<29111> A_IWL<29110> A_IWL<29109> A_IWL<29108> A_IWL<29107> A_IWL<29106> A_IWL<29105> A_IWL<29104> A_IWL<29103> A_IWL<29102> A_IWL<29101> A_IWL<29100> A_IWL<29099> A_IWL<29098> A_IWL<29097> A_IWL<29096> A_IWL<29095> A_IWL<29094> A_IWL<29093> A_IWL<29092> A_IWL<29091> A_IWL<29090> A_IWL<29089> A_IWL<29088> A_IWL<29087> A_IWL<29086> A_IWL<29085> A_IWL<29084> A_IWL<29083> A_IWL<29082> A_IWL<29081> A_IWL<29080> A_IWL<29079> A_IWL<29078> A_IWL<29077> A_IWL<29076> A_IWL<29075> A_IWL<29074> A_IWL<29073> A_IWL<29072> A_IWL<29071> A_IWL<29070> A_IWL<29069> A_IWL<29068> A_IWL<29067> A_IWL<29066> A_IWL<29065> A_IWL<29064> A_IWL<29063> A_IWL<29062> A_IWL<29061> A_IWL<29060> A_IWL<29059> A_IWL<29058> A_IWL<29057> A_IWL<29056> A_IWL<29055> A_IWL<29054> A_IWL<29053> A_IWL<29052> A_IWL<29051> A_IWL<29050> A_IWL<29049> A_IWL<29048> A_IWL<29047> A_IWL<29046> A_IWL<29045> A_IWL<29044> A_IWL<29043> A_IWL<29042> A_IWL<29041> A_IWL<29040> A_IWL<29039> A_IWL<29038> A_IWL<29037> A_IWL<29036> A_IWL<29035> A_IWL<29034> A_IWL<29033> A_IWL<29032> A_IWL<29031> A_IWL<29030> A_IWL<29029> A_IWL<29028> A_IWL<29027> A_IWL<29026> A_IWL<29025> A_IWL<29024> A_IWL<29023> A_IWL<29022> A_IWL<29021> A_IWL<29020> A_IWL<29019> A_IWL<29018> A_IWL<29017> A_IWL<29016> A_IWL<29015> A_IWL<29014> A_IWL<29013> A_IWL<29012> A_IWL<29011> A_IWL<29010> A_IWL<29009> A_IWL<29008> A_IWL<29007> A_IWL<29006> A_IWL<29005> A_IWL<29004> A_IWL<29003> A_IWL<29002> A_IWL<29001> A_IWL<29000> A_IWL<28999> A_IWL<28998> A_IWL<28997> A_IWL<28996> A_IWL<28995> A_IWL<28994> A_IWL<28993> A_IWL<28992> A_IWL<28991> A_IWL<28990> A_IWL<28989> A_IWL<28988> A_IWL<28987> A_IWL<28986> A_IWL<28985> A_IWL<28984> A_IWL<28983> A_IWL<28982> A_IWL<28981> A_IWL<28980> A_IWL<28979> A_IWL<28978> A_IWL<28977> A_IWL<28976> A_IWL<28975> A_IWL<28974> A_IWL<28973> A_IWL<28972> A_IWL<28971> A_IWL<28970> A_IWL<28969> A_IWL<28968> A_IWL<28967> A_IWL<28966> A_IWL<28965> A_IWL<28964> A_IWL<28963> A_IWL<28962> A_IWL<28961> A_IWL<28960> A_IWL<28959> A_IWL<28958> A_IWL<28957> A_IWL<28956> A_IWL<28955> A_IWL<28954> A_IWL<28953> A_IWL<28952> A_IWL<28951> A_IWL<28950> A_IWL<28949> A_IWL<28948> A_IWL<28947> A_IWL<28946> A_IWL<28945> A_IWL<28944> A_IWL<28943> A_IWL<28942> A_IWL<28941> A_IWL<28940> A_IWL<28939> A_IWL<28938> A_IWL<28937> A_IWL<28936> A_IWL<28935> A_IWL<28934> A_IWL<28933> A_IWL<28932> A_IWL<28931> A_IWL<28930> A_IWL<28929> A_IWL<28928> A_IWL<28927> A_IWL<28926> A_IWL<28925> A_IWL<28924> A_IWL<28923> A_IWL<28922> A_IWL<28921> A_IWL<28920> A_IWL<28919> A_IWL<28918> A_IWL<28917> A_IWL<28916> A_IWL<28915> A_IWL<28914> A_IWL<28913> A_IWL<28912> A_IWL<28911> A_IWL<28910> A_IWL<28909> A_IWL<28908> A_IWL<28907> A_IWL<28906> A_IWL<28905> A_IWL<28904> A_IWL<28903> A_IWL<28902> A_IWL<28901> A_IWL<28900> A_IWL<28899> A_IWL<28898> A_IWL<28897> A_IWL<28896> A_IWL<28895> A_IWL<28894> A_IWL<28893> A_IWL<28892> A_IWL<28891> A_IWL<28890> A_IWL<28889> A_IWL<28888> A_IWL<28887> A_IWL<28886> A_IWL<28885> A_IWL<28884> A_IWL<28883> A_IWL<28882> A_IWL<28881> A_IWL<28880> A_IWL<28879> A_IWL<28878> A_IWL<28877> A_IWL<28876> A_IWL<28875> A_IWL<28874> A_IWL<28873> A_IWL<28872> A_IWL<28871> A_IWL<28870> A_IWL<28869> A_IWL<28868> A_IWL<28867> A_IWL<28866> A_IWL<28865> A_IWL<28864> A_IWL<28863> A_IWL<28862> A_IWL<28861> A_IWL<28860> A_IWL<28859> A_IWL<28858> A_IWL<28857> A_IWL<28856> A_IWL<28855> A_IWL<28854> A_IWL<28853> A_IWL<28852> A_IWL<28851> A_IWL<28850> A_IWL<28849> A_IWL<28848> A_IWL<28847> A_IWL<28846> A_IWL<28845> A_IWL<28844> A_IWL<28843> A_IWL<28842> A_IWL<28841> A_IWL<28840> A_IWL<28839> A_IWL<28838> A_IWL<28837> A_IWL<28836> A_IWL<28835> A_IWL<28834> A_IWL<28833> A_IWL<28832> A_IWL<28831> A_IWL<28830> A_IWL<28829> A_IWL<28828> A_IWL<28827> A_IWL<28826> A_IWL<28825> A_IWL<28824> A_IWL<28823> A_IWL<28822> A_IWL<28821> A_IWL<28820> A_IWL<28819> A_IWL<28818> A_IWL<28817> A_IWL<28816> A_IWL<28815> A_IWL<28814> A_IWL<28813> A_IWL<28812> A_IWL<28811> A_IWL<28810> A_IWL<28809> A_IWL<28808> A_IWL<28807> A_IWL<28806> A_IWL<28805> A_IWL<28804> A_IWL<28803> A_IWL<28802> A_IWL<28801> A_IWL<28800> A_IWL<28799> A_IWL<28798> A_IWL<28797> A_IWL<28796> A_IWL<28795> A_IWL<28794> A_IWL<28793> A_IWL<28792> A_IWL<28791> A_IWL<28790> A_IWL<28789> A_IWL<28788> A_IWL<28787> A_IWL<28786> A_IWL<28785> A_IWL<28784> A_IWL<28783> A_IWL<28782> A_IWL<28781> A_IWL<28780> A_IWL<28779> A_IWL<28778> A_IWL<28777> A_IWL<28776> A_IWL<28775> A_IWL<28774> A_IWL<28773> A_IWL<28772> A_IWL<28771> A_IWL<28770> A_IWL<28769> A_IWL<28768> A_IWL<28767> A_IWL<28766> A_IWL<28765> A_IWL<28764> A_IWL<28763> A_IWL<28762> A_IWL<28761> A_IWL<28760> A_IWL<28759> A_IWL<28758> A_IWL<28757> A_IWL<28756> A_IWL<28755> A_IWL<28754> A_IWL<28753> A_IWL<28752> A_IWL<28751> A_IWL<28750> A_IWL<28749> A_IWL<28748> A_IWL<28747> A_IWL<28746> A_IWL<28745> A_IWL<28744> A_IWL<28743> A_IWL<28742> A_IWL<28741> A_IWL<28740> A_IWL<28739> A_IWL<28738> A_IWL<28737> A_IWL<28736> A_IWL<28735> A_IWL<28734> A_IWL<28733> A_IWL<28732> A_IWL<28731> A_IWL<28730> A_IWL<28729> A_IWL<28728> A_IWL<28727> A_IWL<28726> A_IWL<28725> A_IWL<28724> A_IWL<28723> A_IWL<28722> A_IWL<28721> A_IWL<28720> A_IWL<28719> A_IWL<28718> A_IWL<28717> A_IWL<28716> A_IWL<28715> A_IWL<28714> A_IWL<28713> A_IWL<28712> A_IWL<28711> A_IWL<28710> A_IWL<28709> A_IWL<28708> A_IWL<28707> A_IWL<28706> A_IWL<28705> A_IWL<28704> A_IWL<28703> A_IWL<28702> A_IWL<28701> A_IWL<28700> A_IWL<28699> A_IWL<28698> A_IWL<28697> A_IWL<28696> A_IWL<28695> A_IWL<28694> A_IWL<28693> A_IWL<28692> A_IWL<28691> A_IWL<28690> A_IWL<28689> A_IWL<28688> A_IWL<28687> A_IWL<28686> A_IWL<28685> A_IWL<28684> A_IWL<28683> A_IWL<28682> A_IWL<28681> A_IWL<28680> A_IWL<28679> A_IWL<28678> A_IWL<28677> A_IWL<28676> A_IWL<28675> A_IWL<28674> A_IWL<28673> A_IWL<28672> A_IWL<29695> A_IWL<29694> A_IWL<29693> A_IWL<29692> A_IWL<29691> A_IWL<29690> A_IWL<29689> A_IWL<29688> A_IWL<29687> A_IWL<29686> A_IWL<29685> A_IWL<29684> A_IWL<29683> A_IWL<29682> A_IWL<29681> A_IWL<29680> A_IWL<29679> A_IWL<29678> A_IWL<29677> A_IWL<29676> A_IWL<29675> A_IWL<29674> A_IWL<29673> A_IWL<29672> A_IWL<29671> A_IWL<29670> A_IWL<29669> A_IWL<29668> A_IWL<29667> A_IWL<29666> A_IWL<29665> A_IWL<29664> A_IWL<29663> A_IWL<29662> A_IWL<29661> A_IWL<29660> A_IWL<29659> A_IWL<29658> A_IWL<29657> A_IWL<29656> A_IWL<29655> A_IWL<29654> A_IWL<29653> A_IWL<29652> A_IWL<29651> A_IWL<29650> A_IWL<29649> A_IWL<29648> A_IWL<29647> A_IWL<29646> A_IWL<29645> A_IWL<29644> A_IWL<29643> A_IWL<29642> A_IWL<29641> A_IWL<29640> A_IWL<29639> A_IWL<29638> A_IWL<29637> A_IWL<29636> A_IWL<29635> A_IWL<29634> A_IWL<29633> A_IWL<29632> A_IWL<29631> A_IWL<29630> A_IWL<29629> A_IWL<29628> A_IWL<29627> A_IWL<29626> A_IWL<29625> A_IWL<29624> A_IWL<29623> A_IWL<29622> A_IWL<29621> A_IWL<29620> A_IWL<29619> A_IWL<29618> A_IWL<29617> A_IWL<29616> A_IWL<29615> A_IWL<29614> A_IWL<29613> A_IWL<29612> A_IWL<29611> A_IWL<29610> A_IWL<29609> A_IWL<29608> A_IWL<29607> A_IWL<29606> A_IWL<29605> A_IWL<29604> A_IWL<29603> A_IWL<29602> A_IWL<29601> A_IWL<29600> A_IWL<29599> A_IWL<29598> A_IWL<29597> A_IWL<29596> A_IWL<29595> A_IWL<29594> A_IWL<29593> A_IWL<29592> A_IWL<29591> A_IWL<29590> A_IWL<29589> A_IWL<29588> A_IWL<29587> A_IWL<29586> A_IWL<29585> A_IWL<29584> A_IWL<29583> A_IWL<29582> A_IWL<29581> A_IWL<29580> A_IWL<29579> A_IWL<29578> A_IWL<29577> A_IWL<29576> A_IWL<29575> A_IWL<29574> A_IWL<29573> A_IWL<29572> A_IWL<29571> A_IWL<29570> A_IWL<29569> A_IWL<29568> A_IWL<29567> A_IWL<29566> A_IWL<29565> A_IWL<29564> A_IWL<29563> A_IWL<29562> A_IWL<29561> A_IWL<29560> A_IWL<29559> A_IWL<29558> A_IWL<29557> A_IWL<29556> A_IWL<29555> A_IWL<29554> A_IWL<29553> A_IWL<29552> A_IWL<29551> A_IWL<29550> A_IWL<29549> A_IWL<29548> A_IWL<29547> A_IWL<29546> A_IWL<29545> A_IWL<29544> A_IWL<29543> A_IWL<29542> A_IWL<29541> A_IWL<29540> A_IWL<29539> A_IWL<29538> A_IWL<29537> A_IWL<29536> A_IWL<29535> A_IWL<29534> A_IWL<29533> A_IWL<29532> A_IWL<29531> A_IWL<29530> A_IWL<29529> A_IWL<29528> A_IWL<29527> A_IWL<29526> A_IWL<29525> A_IWL<29524> A_IWL<29523> A_IWL<29522> A_IWL<29521> A_IWL<29520> A_IWL<29519> A_IWL<29518> A_IWL<29517> A_IWL<29516> A_IWL<29515> A_IWL<29514> A_IWL<29513> A_IWL<29512> A_IWL<29511> A_IWL<29510> A_IWL<29509> A_IWL<29508> A_IWL<29507> A_IWL<29506> A_IWL<29505> A_IWL<29504> A_IWL<29503> A_IWL<29502> A_IWL<29501> A_IWL<29500> A_IWL<29499> A_IWL<29498> A_IWL<29497> A_IWL<29496> A_IWL<29495> A_IWL<29494> A_IWL<29493> A_IWL<29492> A_IWL<29491> A_IWL<29490> A_IWL<29489> A_IWL<29488> A_IWL<29487> A_IWL<29486> A_IWL<29485> A_IWL<29484> A_IWL<29483> A_IWL<29482> A_IWL<29481> A_IWL<29480> A_IWL<29479> A_IWL<29478> A_IWL<29477> A_IWL<29476> A_IWL<29475> A_IWL<29474> A_IWL<29473> A_IWL<29472> A_IWL<29471> A_IWL<29470> A_IWL<29469> A_IWL<29468> A_IWL<29467> A_IWL<29466> A_IWL<29465> A_IWL<29464> A_IWL<29463> A_IWL<29462> A_IWL<29461> A_IWL<29460> A_IWL<29459> A_IWL<29458> A_IWL<29457> A_IWL<29456> A_IWL<29455> A_IWL<29454> A_IWL<29453> A_IWL<29452> A_IWL<29451> A_IWL<29450> A_IWL<29449> A_IWL<29448> A_IWL<29447> A_IWL<29446> A_IWL<29445> A_IWL<29444> A_IWL<29443> A_IWL<29442> A_IWL<29441> A_IWL<29440> A_IWL<29439> A_IWL<29438> A_IWL<29437> A_IWL<29436> A_IWL<29435> A_IWL<29434> A_IWL<29433> A_IWL<29432> A_IWL<29431> A_IWL<29430> A_IWL<29429> A_IWL<29428> A_IWL<29427> A_IWL<29426> A_IWL<29425> A_IWL<29424> A_IWL<29423> A_IWL<29422> A_IWL<29421> A_IWL<29420> A_IWL<29419> A_IWL<29418> A_IWL<29417> A_IWL<29416> A_IWL<29415> A_IWL<29414> A_IWL<29413> A_IWL<29412> A_IWL<29411> A_IWL<29410> A_IWL<29409> A_IWL<29408> A_IWL<29407> A_IWL<29406> A_IWL<29405> A_IWL<29404> A_IWL<29403> A_IWL<29402> A_IWL<29401> A_IWL<29400> A_IWL<29399> A_IWL<29398> A_IWL<29397> A_IWL<29396> A_IWL<29395> A_IWL<29394> A_IWL<29393> A_IWL<29392> A_IWL<29391> A_IWL<29390> A_IWL<29389> A_IWL<29388> A_IWL<29387> A_IWL<29386> A_IWL<29385> A_IWL<29384> A_IWL<29383> A_IWL<29382> A_IWL<29381> A_IWL<29380> A_IWL<29379> A_IWL<29378> A_IWL<29377> A_IWL<29376> A_IWL<29375> A_IWL<29374> A_IWL<29373> A_IWL<29372> A_IWL<29371> A_IWL<29370> A_IWL<29369> A_IWL<29368> A_IWL<29367> A_IWL<29366> A_IWL<29365> A_IWL<29364> A_IWL<29363> A_IWL<29362> A_IWL<29361> A_IWL<29360> A_IWL<29359> A_IWL<29358> A_IWL<29357> A_IWL<29356> A_IWL<29355> A_IWL<29354> A_IWL<29353> A_IWL<29352> A_IWL<29351> A_IWL<29350> A_IWL<29349> A_IWL<29348> A_IWL<29347> A_IWL<29346> A_IWL<29345> A_IWL<29344> A_IWL<29343> A_IWL<29342> A_IWL<29341> A_IWL<29340> A_IWL<29339> A_IWL<29338> A_IWL<29337> A_IWL<29336> A_IWL<29335> A_IWL<29334> A_IWL<29333> A_IWL<29332> A_IWL<29331> A_IWL<29330> A_IWL<29329> A_IWL<29328> A_IWL<29327> A_IWL<29326> A_IWL<29325> A_IWL<29324> A_IWL<29323> A_IWL<29322> A_IWL<29321> A_IWL<29320> A_IWL<29319> A_IWL<29318> A_IWL<29317> A_IWL<29316> A_IWL<29315> A_IWL<29314> A_IWL<29313> A_IWL<29312> A_IWL<29311> A_IWL<29310> A_IWL<29309> A_IWL<29308> A_IWL<29307> A_IWL<29306> A_IWL<29305> A_IWL<29304> A_IWL<29303> A_IWL<29302> A_IWL<29301> A_IWL<29300> A_IWL<29299> A_IWL<29298> A_IWL<29297> A_IWL<29296> A_IWL<29295> A_IWL<29294> A_IWL<29293> A_IWL<29292> A_IWL<29291> A_IWL<29290> A_IWL<29289> A_IWL<29288> A_IWL<29287> A_IWL<29286> A_IWL<29285> A_IWL<29284> A_IWL<29283> A_IWL<29282> A_IWL<29281> A_IWL<29280> A_IWL<29279> A_IWL<29278> A_IWL<29277> A_IWL<29276> A_IWL<29275> A_IWL<29274> A_IWL<29273> A_IWL<29272> A_IWL<29271> A_IWL<29270> A_IWL<29269> A_IWL<29268> A_IWL<29267> A_IWL<29266> A_IWL<29265> A_IWL<29264> A_IWL<29263> A_IWL<29262> A_IWL<29261> A_IWL<29260> A_IWL<29259> A_IWL<29258> A_IWL<29257> A_IWL<29256> A_IWL<29255> A_IWL<29254> A_IWL<29253> A_IWL<29252> A_IWL<29251> A_IWL<29250> A_IWL<29249> A_IWL<29248> A_IWL<29247> A_IWL<29246> A_IWL<29245> A_IWL<29244> A_IWL<29243> A_IWL<29242> A_IWL<29241> A_IWL<29240> A_IWL<29239> A_IWL<29238> A_IWL<29237> A_IWL<29236> A_IWL<29235> A_IWL<29234> A_IWL<29233> A_IWL<29232> A_IWL<29231> A_IWL<29230> A_IWL<29229> A_IWL<29228> A_IWL<29227> A_IWL<29226> A_IWL<29225> A_IWL<29224> A_IWL<29223> A_IWL<29222> A_IWL<29221> A_IWL<29220> A_IWL<29219> A_IWL<29218> A_IWL<29217> A_IWL<29216> A_IWL<29215> A_IWL<29214> A_IWL<29213> A_IWL<29212> A_IWL<29211> A_IWL<29210> A_IWL<29209> A_IWL<29208> A_IWL<29207> A_IWL<29206> A_IWL<29205> A_IWL<29204> A_IWL<29203> A_IWL<29202> A_IWL<29201> A_IWL<29200> A_IWL<29199> A_IWL<29198> A_IWL<29197> A_IWL<29196> A_IWL<29195> A_IWL<29194> A_IWL<29193> A_IWL<29192> A_IWL<29191> A_IWL<29190> A_IWL<29189> A_IWL<29188> A_IWL<29187> A_IWL<29186> A_IWL<29185> A_IWL<29184> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<56> A_BLC<113> A_BLC<112> A_BLC_TOP<113> A_BLC_TOP<112> A_BLT<113> A_BLT<112> A_BLT_TOP<113> A_BLT_TOP<112> A_IWL<28671> A_IWL<28670> A_IWL<28669> A_IWL<28668> A_IWL<28667> A_IWL<28666> A_IWL<28665> A_IWL<28664> A_IWL<28663> A_IWL<28662> A_IWL<28661> A_IWL<28660> A_IWL<28659> A_IWL<28658> A_IWL<28657> A_IWL<28656> A_IWL<28655> A_IWL<28654> A_IWL<28653> A_IWL<28652> A_IWL<28651> A_IWL<28650> A_IWL<28649> A_IWL<28648> A_IWL<28647> A_IWL<28646> A_IWL<28645> A_IWL<28644> A_IWL<28643> A_IWL<28642> A_IWL<28641> A_IWL<28640> A_IWL<28639> A_IWL<28638> A_IWL<28637> A_IWL<28636> A_IWL<28635> A_IWL<28634> A_IWL<28633> A_IWL<28632> A_IWL<28631> A_IWL<28630> A_IWL<28629> A_IWL<28628> A_IWL<28627> A_IWL<28626> A_IWL<28625> A_IWL<28624> A_IWL<28623> A_IWL<28622> A_IWL<28621> A_IWL<28620> A_IWL<28619> A_IWL<28618> A_IWL<28617> A_IWL<28616> A_IWL<28615> A_IWL<28614> A_IWL<28613> A_IWL<28612> A_IWL<28611> A_IWL<28610> A_IWL<28609> A_IWL<28608> A_IWL<28607> A_IWL<28606> A_IWL<28605> A_IWL<28604> A_IWL<28603> A_IWL<28602> A_IWL<28601> A_IWL<28600> A_IWL<28599> A_IWL<28598> A_IWL<28597> A_IWL<28596> A_IWL<28595> A_IWL<28594> A_IWL<28593> A_IWL<28592> A_IWL<28591> A_IWL<28590> A_IWL<28589> A_IWL<28588> A_IWL<28587> A_IWL<28586> A_IWL<28585> A_IWL<28584> A_IWL<28583> A_IWL<28582> A_IWL<28581> A_IWL<28580> A_IWL<28579> A_IWL<28578> A_IWL<28577> A_IWL<28576> A_IWL<28575> A_IWL<28574> A_IWL<28573> A_IWL<28572> A_IWL<28571> A_IWL<28570> A_IWL<28569> A_IWL<28568> A_IWL<28567> A_IWL<28566> A_IWL<28565> A_IWL<28564> A_IWL<28563> A_IWL<28562> A_IWL<28561> A_IWL<28560> A_IWL<28559> A_IWL<28558> A_IWL<28557> A_IWL<28556> A_IWL<28555> A_IWL<28554> A_IWL<28553> A_IWL<28552> A_IWL<28551> A_IWL<28550> A_IWL<28549> A_IWL<28548> A_IWL<28547> A_IWL<28546> A_IWL<28545> A_IWL<28544> A_IWL<28543> A_IWL<28542> A_IWL<28541> A_IWL<28540> A_IWL<28539> A_IWL<28538> A_IWL<28537> A_IWL<28536> A_IWL<28535> A_IWL<28534> A_IWL<28533> A_IWL<28532> A_IWL<28531> A_IWL<28530> A_IWL<28529> A_IWL<28528> A_IWL<28527> A_IWL<28526> A_IWL<28525> A_IWL<28524> A_IWL<28523> A_IWL<28522> A_IWL<28521> A_IWL<28520> A_IWL<28519> A_IWL<28518> A_IWL<28517> A_IWL<28516> A_IWL<28515> A_IWL<28514> A_IWL<28513> A_IWL<28512> A_IWL<28511> A_IWL<28510> A_IWL<28509> A_IWL<28508> A_IWL<28507> A_IWL<28506> A_IWL<28505> A_IWL<28504> A_IWL<28503> A_IWL<28502> A_IWL<28501> A_IWL<28500> A_IWL<28499> A_IWL<28498> A_IWL<28497> A_IWL<28496> A_IWL<28495> A_IWL<28494> A_IWL<28493> A_IWL<28492> A_IWL<28491> A_IWL<28490> A_IWL<28489> A_IWL<28488> A_IWL<28487> A_IWL<28486> A_IWL<28485> A_IWL<28484> A_IWL<28483> A_IWL<28482> A_IWL<28481> A_IWL<28480> A_IWL<28479> A_IWL<28478> A_IWL<28477> A_IWL<28476> A_IWL<28475> A_IWL<28474> A_IWL<28473> A_IWL<28472> A_IWL<28471> A_IWL<28470> A_IWL<28469> A_IWL<28468> A_IWL<28467> A_IWL<28466> A_IWL<28465> A_IWL<28464> A_IWL<28463> A_IWL<28462> A_IWL<28461> A_IWL<28460> A_IWL<28459> A_IWL<28458> A_IWL<28457> A_IWL<28456> A_IWL<28455> A_IWL<28454> A_IWL<28453> A_IWL<28452> A_IWL<28451> A_IWL<28450> A_IWL<28449> A_IWL<28448> A_IWL<28447> A_IWL<28446> A_IWL<28445> A_IWL<28444> A_IWL<28443> A_IWL<28442> A_IWL<28441> A_IWL<28440> A_IWL<28439> A_IWL<28438> A_IWL<28437> A_IWL<28436> A_IWL<28435> A_IWL<28434> A_IWL<28433> A_IWL<28432> A_IWL<28431> A_IWL<28430> A_IWL<28429> A_IWL<28428> A_IWL<28427> A_IWL<28426> A_IWL<28425> A_IWL<28424> A_IWL<28423> A_IWL<28422> A_IWL<28421> A_IWL<28420> A_IWL<28419> A_IWL<28418> A_IWL<28417> A_IWL<28416> A_IWL<28415> A_IWL<28414> A_IWL<28413> A_IWL<28412> A_IWL<28411> A_IWL<28410> A_IWL<28409> A_IWL<28408> A_IWL<28407> A_IWL<28406> A_IWL<28405> A_IWL<28404> A_IWL<28403> A_IWL<28402> A_IWL<28401> A_IWL<28400> A_IWL<28399> A_IWL<28398> A_IWL<28397> A_IWL<28396> A_IWL<28395> A_IWL<28394> A_IWL<28393> A_IWL<28392> A_IWL<28391> A_IWL<28390> A_IWL<28389> A_IWL<28388> A_IWL<28387> A_IWL<28386> A_IWL<28385> A_IWL<28384> A_IWL<28383> A_IWL<28382> A_IWL<28381> A_IWL<28380> A_IWL<28379> A_IWL<28378> A_IWL<28377> A_IWL<28376> A_IWL<28375> A_IWL<28374> A_IWL<28373> A_IWL<28372> A_IWL<28371> A_IWL<28370> A_IWL<28369> A_IWL<28368> A_IWL<28367> A_IWL<28366> A_IWL<28365> A_IWL<28364> A_IWL<28363> A_IWL<28362> A_IWL<28361> A_IWL<28360> A_IWL<28359> A_IWL<28358> A_IWL<28357> A_IWL<28356> A_IWL<28355> A_IWL<28354> A_IWL<28353> A_IWL<28352> A_IWL<28351> A_IWL<28350> A_IWL<28349> A_IWL<28348> A_IWL<28347> A_IWL<28346> A_IWL<28345> A_IWL<28344> A_IWL<28343> A_IWL<28342> A_IWL<28341> A_IWL<28340> A_IWL<28339> A_IWL<28338> A_IWL<28337> A_IWL<28336> A_IWL<28335> A_IWL<28334> A_IWL<28333> A_IWL<28332> A_IWL<28331> A_IWL<28330> A_IWL<28329> A_IWL<28328> A_IWL<28327> A_IWL<28326> A_IWL<28325> A_IWL<28324> A_IWL<28323> A_IWL<28322> A_IWL<28321> A_IWL<28320> A_IWL<28319> A_IWL<28318> A_IWL<28317> A_IWL<28316> A_IWL<28315> A_IWL<28314> A_IWL<28313> A_IWL<28312> A_IWL<28311> A_IWL<28310> A_IWL<28309> A_IWL<28308> A_IWL<28307> A_IWL<28306> A_IWL<28305> A_IWL<28304> A_IWL<28303> A_IWL<28302> A_IWL<28301> A_IWL<28300> A_IWL<28299> A_IWL<28298> A_IWL<28297> A_IWL<28296> A_IWL<28295> A_IWL<28294> A_IWL<28293> A_IWL<28292> A_IWL<28291> A_IWL<28290> A_IWL<28289> A_IWL<28288> A_IWL<28287> A_IWL<28286> A_IWL<28285> A_IWL<28284> A_IWL<28283> A_IWL<28282> A_IWL<28281> A_IWL<28280> A_IWL<28279> A_IWL<28278> A_IWL<28277> A_IWL<28276> A_IWL<28275> A_IWL<28274> A_IWL<28273> A_IWL<28272> A_IWL<28271> A_IWL<28270> A_IWL<28269> A_IWL<28268> A_IWL<28267> A_IWL<28266> A_IWL<28265> A_IWL<28264> A_IWL<28263> A_IWL<28262> A_IWL<28261> A_IWL<28260> A_IWL<28259> A_IWL<28258> A_IWL<28257> A_IWL<28256> A_IWL<28255> A_IWL<28254> A_IWL<28253> A_IWL<28252> A_IWL<28251> A_IWL<28250> A_IWL<28249> A_IWL<28248> A_IWL<28247> A_IWL<28246> A_IWL<28245> A_IWL<28244> A_IWL<28243> A_IWL<28242> A_IWL<28241> A_IWL<28240> A_IWL<28239> A_IWL<28238> A_IWL<28237> A_IWL<28236> A_IWL<28235> A_IWL<28234> A_IWL<28233> A_IWL<28232> A_IWL<28231> A_IWL<28230> A_IWL<28229> A_IWL<28228> A_IWL<28227> A_IWL<28226> A_IWL<28225> A_IWL<28224> A_IWL<28223> A_IWL<28222> A_IWL<28221> A_IWL<28220> A_IWL<28219> A_IWL<28218> A_IWL<28217> A_IWL<28216> A_IWL<28215> A_IWL<28214> A_IWL<28213> A_IWL<28212> A_IWL<28211> A_IWL<28210> A_IWL<28209> A_IWL<28208> A_IWL<28207> A_IWL<28206> A_IWL<28205> A_IWL<28204> A_IWL<28203> A_IWL<28202> A_IWL<28201> A_IWL<28200> A_IWL<28199> A_IWL<28198> A_IWL<28197> A_IWL<28196> A_IWL<28195> A_IWL<28194> A_IWL<28193> A_IWL<28192> A_IWL<28191> A_IWL<28190> A_IWL<28189> A_IWL<28188> A_IWL<28187> A_IWL<28186> A_IWL<28185> A_IWL<28184> A_IWL<28183> A_IWL<28182> A_IWL<28181> A_IWL<28180> A_IWL<28179> A_IWL<28178> A_IWL<28177> A_IWL<28176> A_IWL<28175> A_IWL<28174> A_IWL<28173> A_IWL<28172> A_IWL<28171> A_IWL<28170> A_IWL<28169> A_IWL<28168> A_IWL<28167> A_IWL<28166> A_IWL<28165> A_IWL<28164> A_IWL<28163> A_IWL<28162> A_IWL<28161> A_IWL<28160> A_IWL<29183> A_IWL<29182> A_IWL<29181> A_IWL<29180> A_IWL<29179> A_IWL<29178> A_IWL<29177> A_IWL<29176> A_IWL<29175> A_IWL<29174> A_IWL<29173> A_IWL<29172> A_IWL<29171> A_IWL<29170> A_IWL<29169> A_IWL<29168> A_IWL<29167> A_IWL<29166> A_IWL<29165> A_IWL<29164> A_IWL<29163> A_IWL<29162> A_IWL<29161> A_IWL<29160> A_IWL<29159> A_IWL<29158> A_IWL<29157> A_IWL<29156> A_IWL<29155> A_IWL<29154> A_IWL<29153> A_IWL<29152> A_IWL<29151> A_IWL<29150> A_IWL<29149> A_IWL<29148> A_IWL<29147> A_IWL<29146> A_IWL<29145> A_IWL<29144> A_IWL<29143> A_IWL<29142> A_IWL<29141> A_IWL<29140> A_IWL<29139> A_IWL<29138> A_IWL<29137> A_IWL<29136> A_IWL<29135> A_IWL<29134> A_IWL<29133> A_IWL<29132> A_IWL<29131> A_IWL<29130> A_IWL<29129> A_IWL<29128> A_IWL<29127> A_IWL<29126> A_IWL<29125> A_IWL<29124> A_IWL<29123> A_IWL<29122> A_IWL<29121> A_IWL<29120> A_IWL<29119> A_IWL<29118> A_IWL<29117> A_IWL<29116> A_IWL<29115> A_IWL<29114> A_IWL<29113> A_IWL<29112> A_IWL<29111> A_IWL<29110> A_IWL<29109> A_IWL<29108> A_IWL<29107> A_IWL<29106> A_IWL<29105> A_IWL<29104> A_IWL<29103> A_IWL<29102> A_IWL<29101> A_IWL<29100> A_IWL<29099> A_IWL<29098> A_IWL<29097> A_IWL<29096> A_IWL<29095> A_IWL<29094> A_IWL<29093> A_IWL<29092> A_IWL<29091> A_IWL<29090> A_IWL<29089> A_IWL<29088> A_IWL<29087> A_IWL<29086> A_IWL<29085> A_IWL<29084> A_IWL<29083> A_IWL<29082> A_IWL<29081> A_IWL<29080> A_IWL<29079> A_IWL<29078> A_IWL<29077> A_IWL<29076> A_IWL<29075> A_IWL<29074> A_IWL<29073> A_IWL<29072> A_IWL<29071> A_IWL<29070> A_IWL<29069> A_IWL<29068> A_IWL<29067> A_IWL<29066> A_IWL<29065> A_IWL<29064> A_IWL<29063> A_IWL<29062> A_IWL<29061> A_IWL<29060> A_IWL<29059> A_IWL<29058> A_IWL<29057> A_IWL<29056> A_IWL<29055> A_IWL<29054> A_IWL<29053> A_IWL<29052> A_IWL<29051> A_IWL<29050> A_IWL<29049> A_IWL<29048> A_IWL<29047> A_IWL<29046> A_IWL<29045> A_IWL<29044> A_IWL<29043> A_IWL<29042> A_IWL<29041> A_IWL<29040> A_IWL<29039> A_IWL<29038> A_IWL<29037> A_IWL<29036> A_IWL<29035> A_IWL<29034> A_IWL<29033> A_IWL<29032> A_IWL<29031> A_IWL<29030> A_IWL<29029> A_IWL<29028> A_IWL<29027> A_IWL<29026> A_IWL<29025> A_IWL<29024> A_IWL<29023> A_IWL<29022> A_IWL<29021> A_IWL<29020> A_IWL<29019> A_IWL<29018> A_IWL<29017> A_IWL<29016> A_IWL<29015> A_IWL<29014> A_IWL<29013> A_IWL<29012> A_IWL<29011> A_IWL<29010> A_IWL<29009> A_IWL<29008> A_IWL<29007> A_IWL<29006> A_IWL<29005> A_IWL<29004> A_IWL<29003> A_IWL<29002> A_IWL<29001> A_IWL<29000> A_IWL<28999> A_IWL<28998> A_IWL<28997> A_IWL<28996> A_IWL<28995> A_IWL<28994> A_IWL<28993> A_IWL<28992> A_IWL<28991> A_IWL<28990> A_IWL<28989> A_IWL<28988> A_IWL<28987> A_IWL<28986> A_IWL<28985> A_IWL<28984> A_IWL<28983> A_IWL<28982> A_IWL<28981> A_IWL<28980> A_IWL<28979> A_IWL<28978> A_IWL<28977> A_IWL<28976> A_IWL<28975> A_IWL<28974> A_IWL<28973> A_IWL<28972> A_IWL<28971> A_IWL<28970> A_IWL<28969> A_IWL<28968> A_IWL<28967> A_IWL<28966> A_IWL<28965> A_IWL<28964> A_IWL<28963> A_IWL<28962> A_IWL<28961> A_IWL<28960> A_IWL<28959> A_IWL<28958> A_IWL<28957> A_IWL<28956> A_IWL<28955> A_IWL<28954> A_IWL<28953> A_IWL<28952> A_IWL<28951> A_IWL<28950> A_IWL<28949> A_IWL<28948> A_IWL<28947> A_IWL<28946> A_IWL<28945> A_IWL<28944> A_IWL<28943> A_IWL<28942> A_IWL<28941> A_IWL<28940> A_IWL<28939> A_IWL<28938> A_IWL<28937> A_IWL<28936> A_IWL<28935> A_IWL<28934> A_IWL<28933> A_IWL<28932> A_IWL<28931> A_IWL<28930> A_IWL<28929> A_IWL<28928> A_IWL<28927> A_IWL<28926> A_IWL<28925> A_IWL<28924> A_IWL<28923> A_IWL<28922> A_IWL<28921> A_IWL<28920> A_IWL<28919> A_IWL<28918> A_IWL<28917> A_IWL<28916> A_IWL<28915> A_IWL<28914> A_IWL<28913> A_IWL<28912> A_IWL<28911> A_IWL<28910> A_IWL<28909> A_IWL<28908> A_IWL<28907> A_IWL<28906> A_IWL<28905> A_IWL<28904> A_IWL<28903> A_IWL<28902> A_IWL<28901> A_IWL<28900> A_IWL<28899> A_IWL<28898> A_IWL<28897> A_IWL<28896> A_IWL<28895> A_IWL<28894> A_IWL<28893> A_IWL<28892> A_IWL<28891> A_IWL<28890> A_IWL<28889> A_IWL<28888> A_IWL<28887> A_IWL<28886> A_IWL<28885> A_IWL<28884> A_IWL<28883> A_IWL<28882> A_IWL<28881> A_IWL<28880> A_IWL<28879> A_IWL<28878> A_IWL<28877> A_IWL<28876> A_IWL<28875> A_IWL<28874> A_IWL<28873> A_IWL<28872> A_IWL<28871> A_IWL<28870> A_IWL<28869> A_IWL<28868> A_IWL<28867> A_IWL<28866> A_IWL<28865> A_IWL<28864> A_IWL<28863> A_IWL<28862> A_IWL<28861> A_IWL<28860> A_IWL<28859> A_IWL<28858> A_IWL<28857> A_IWL<28856> A_IWL<28855> A_IWL<28854> A_IWL<28853> A_IWL<28852> A_IWL<28851> A_IWL<28850> A_IWL<28849> A_IWL<28848> A_IWL<28847> A_IWL<28846> A_IWL<28845> A_IWL<28844> A_IWL<28843> A_IWL<28842> A_IWL<28841> A_IWL<28840> A_IWL<28839> A_IWL<28838> A_IWL<28837> A_IWL<28836> A_IWL<28835> A_IWL<28834> A_IWL<28833> A_IWL<28832> A_IWL<28831> A_IWL<28830> A_IWL<28829> A_IWL<28828> A_IWL<28827> A_IWL<28826> A_IWL<28825> A_IWL<28824> A_IWL<28823> A_IWL<28822> A_IWL<28821> A_IWL<28820> A_IWL<28819> A_IWL<28818> A_IWL<28817> A_IWL<28816> A_IWL<28815> A_IWL<28814> A_IWL<28813> A_IWL<28812> A_IWL<28811> A_IWL<28810> A_IWL<28809> A_IWL<28808> A_IWL<28807> A_IWL<28806> A_IWL<28805> A_IWL<28804> A_IWL<28803> A_IWL<28802> A_IWL<28801> A_IWL<28800> A_IWL<28799> A_IWL<28798> A_IWL<28797> A_IWL<28796> A_IWL<28795> A_IWL<28794> A_IWL<28793> A_IWL<28792> A_IWL<28791> A_IWL<28790> A_IWL<28789> A_IWL<28788> A_IWL<28787> A_IWL<28786> A_IWL<28785> A_IWL<28784> A_IWL<28783> A_IWL<28782> A_IWL<28781> A_IWL<28780> A_IWL<28779> A_IWL<28778> A_IWL<28777> A_IWL<28776> A_IWL<28775> A_IWL<28774> A_IWL<28773> A_IWL<28772> A_IWL<28771> A_IWL<28770> A_IWL<28769> A_IWL<28768> A_IWL<28767> A_IWL<28766> A_IWL<28765> A_IWL<28764> A_IWL<28763> A_IWL<28762> A_IWL<28761> A_IWL<28760> A_IWL<28759> A_IWL<28758> A_IWL<28757> A_IWL<28756> A_IWL<28755> A_IWL<28754> A_IWL<28753> A_IWL<28752> A_IWL<28751> A_IWL<28750> A_IWL<28749> A_IWL<28748> A_IWL<28747> A_IWL<28746> A_IWL<28745> A_IWL<28744> A_IWL<28743> A_IWL<28742> A_IWL<28741> A_IWL<28740> A_IWL<28739> A_IWL<28738> A_IWL<28737> A_IWL<28736> A_IWL<28735> A_IWL<28734> A_IWL<28733> A_IWL<28732> A_IWL<28731> A_IWL<28730> A_IWL<28729> A_IWL<28728> A_IWL<28727> A_IWL<28726> A_IWL<28725> A_IWL<28724> A_IWL<28723> A_IWL<28722> A_IWL<28721> A_IWL<28720> A_IWL<28719> A_IWL<28718> A_IWL<28717> A_IWL<28716> A_IWL<28715> A_IWL<28714> A_IWL<28713> A_IWL<28712> A_IWL<28711> A_IWL<28710> A_IWL<28709> A_IWL<28708> A_IWL<28707> A_IWL<28706> A_IWL<28705> A_IWL<28704> A_IWL<28703> A_IWL<28702> A_IWL<28701> A_IWL<28700> A_IWL<28699> A_IWL<28698> A_IWL<28697> A_IWL<28696> A_IWL<28695> A_IWL<28694> A_IWL<28693> A_IWL<28692> A_IWL<28691> A_IWL<28690> A_IWL<28689> A_IWL<28688> A_IWL<28687> A_IWL<28686> A_IWL<28685> A_IWL<28684> A_IWL<28683> A_IWL<28682> A_IWL<28681> A_IWL<28680> A_IWL<28679> A_IWL<28678> A_IWL<28677> A_IWL<28676> A_IWL<28675> A_IWL<28674> A_IWL<28673> A_IWL<28672> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<55> A_BLC<111> A_BLC<110> A_BLC_TOP<111> A_BLC_TOP<110> A_BLT<111> A_BLT<110> A_BLT_TOP<111> A_BLT_TOP<110> A_IWL<28159> A_IWL<28158> A_IWL<28157> A_IWL<28156> A_IWL<28155> A_IWL<28154> A_IWL<28153> A_IWL<28152> A_IWL<28151> A_IWL<28150> A_IWL<28149> A_IWL<28148> A_IWL<28147> A_IWL<28146> A_IWL<28145> A_IWL<28144> A_IWL<28143> A_IWL<28142> A_IWL<28141> A_IWL<28140> A_IWL<28139> A_IWL<28138> A_IWL<28137> A_IWL<28136> A_IWL<28135> A_IWL<28134> A_IWL<28133> A_IWL<28132> A_IWL<28131> A_IWL<28130> A_IWL<28129> A_IWL<28128> A_IWL<28127> A_IWL<28126> A_IWL<28125> A_IWL<28124> A_IWL<28123> A_IWL<28122> A_IWL<28121> A_IWL<28120> A_IWL<28119> A_IWL<28118> A_IWL<28117> A_IWL<28116> A_IWL<28115> A_IWL<28114> A_IWL<28113> A_IWL<28112> A_IWL<28111> A_IWL<28110> A_IWL<28109> A_IWL<28108> A_IWL<28107> A_IWL<28106> A_IWL<28105> A_IWL<28104> A_IWL<28103> A_IWL<28102> A_IWL<28101> A_IWL<28100> A_IWL<28099> A_IWL<28098> A_IWL<28097> A_IWL<28096> A_IWL<28095> A_IWL<28094> A_IWL<28093> A_IWL<28092> A_IWL<28091> A_IWL<28090> A_IWL<28089> A_IWL<28088> A_IWL<28087> A_IWL<28086> A_IWL<28085> A_IWL<28084> A_IWL<28083> A_IWL<28082> A_IWL<28081> A_IWL<28080> A_IWL<28079> A_IWL<28078> A_IWL<28077> A_IWL<28076> A_IWL<28075> A_IWL<28074> A_IWL<28073> A_IWL<28072> A_IWL<28071> A_IWL<28070> A_IWL<28069> A_IWL<28068> A_IWL<28067> A_IWL<28066> A_IWL<28065> A_IWL<28064> A_IWL<28063> A_IWL<28062> A_IWL<28061> A_IWL<28060> A_IWL<28059> A_IWL<28058> A_IWL<28057> A_IWL<28056> A_IWL<28055> A_IWL<28054> A_IWL<28053> A_IWL<28052> A_IWL<28051> A_IWL<28050> A_IWL<28049> A_IWL<28048> A_IWL<28047> A_IWL<28046> A_IWL<28045> A_IWL<28044> A_IWL<28043> A_IWL<28042> A_IWL<28041> A_IWL<28040> A_IWL<28039> A_IWL<28038> A_IWL<28037> A_IWL<28036> A_IWL<28035> A_IWL<28034> A_IWL<28033> A_IWL<28032> A_IWL<28031> A_IWL<28030> A_IWL<28029> A_IWL<28028> A_IWL<28027> A_IWL<28026> A_IWL<28025> A_IWL<28024> A_IWL<28023> A_IWL<28022> A_IWL<28021> A_IWL<28020> A_IWL<28019> A_IWL<28018> A_IWL<28017> A_IWL<28016> A_IWL<28015> A_IWL<28014> A_IWL<28013> A_IWL<28012> A_IWL<28011> A_IWL<28010> A_IWL<28009> A_IWL<28008> A_IWL<28007> A_IWL<28006> A_IWL<28005> A_IWL<28004> A_IWL<28003> A_IWL<28002> A_IWL<28001> A_IWL<28000> A_IWL<27999> A_IWL<27998> A_IWL<27997> A_IWL<27996> A_IWL<27995> A_IWL<27994> A_IWL<27993> A_IWL<27992> A_IWL<27991> A_IWL<27990> A_IWL<27989> A_IWL<27988> A_IWL<27987> A_IWL<27986> A_IWL<27985> A_IWL<27984> A_IWL<27983> A_IWL<27982> A_IWL<27981> A_IWL<27980> A_IWL<27979> A_IWL<27978> A_IWL<27977> A_IWL<27976> A_IWL<27975> A_IWL<27974> A_IWL<27973> A_IWL<27972> A_IWL<27971> A_IWL<27970> A_IWL<27969> A_IWL<27968> A_IWL<27967> A_IWL<27966> A_IWL<27965> A_IWL<27964> A_IWL<27963> A_IWL<27962> A_IWL<27961> A_IWL<27960> A_IWL<27959> A_IWL<27958> A_IWL<27957> A_IWL<27956> A_IWL<27955> A_IWL<27954> A_IWL<27953> A_IWL<27952> A_IWL<27951> A_IWL<27950> A_IWL<27949> A_IWL<27948> A_IWL<27947> A_IWL<27946> A_IWL<27945> A_IWL<27944> A_IWL<27943> A_IWL<27942> A_IWL<27941> A_IWL<27940> A_IWL<27939> A_IWL<27938> A_IWL<27937> A_IWL<27936> A_IWL<27935> A_IWL<27934> A_IWL<27933> A_IWL<27932> A_IWL<27931> A_IWL<27930> A_IWL<27929> A_IWL<27928> A_IWL<27927> A_IWL<27926> A_IWL<27925> A_IWL<27924> A_IWL<27923> A_IWL<27922> A_IWL<27921> A_IWL<27920> A_IWL<27919> A_IWL<27918> A_IWL<27917> A_IWL<27916> A_IWL<27915> A_IWL<27914> A_IWL<27913> A_IWL<27912> A_IWL<27911> A_IWL<27910> A_IWL<27909> A_IWL<27908> A_IWL<27907> A_IWL<27906> A_IWL<27905> A_IWL<27904> A_IWL<27903> A_IWL<27902> A_IWL<27901> A_IWL<27900> A_IWL<27899> A_IWL<27898> A_IWL<27897> A_IWL<27896> A_IWL<27895> A_IWL<27894> A_IWL<27893> A_IWL<27892> A_IWL<27891> A_IWL<27890> A_IWL<27889> A_IWL<27888> A_IWL<27887> A_IWL<27886> A_IWL<27885> A_IWL<27884> A_IWL<27883> A_IWL<27882> A_IWL<27881> A_IWL<27880> A_IWL<27879> A_IWL<27878> A_IWL<27877> A_IWL<27876> A_IWL<27875> A_IWL<27874> A_IWL<27873> A_IWL<27872> A_IWL<27871> A_IWL<27870> A_IWL<27869> A_IWL<27868> A_IWL<27867> A_IWL<27866> A_IWL<27865> A_IWL<27864> A_IWL<27863> A_IWL<27862> A_IWL<27861> A_IWL<27860> A_IWL<27859> A_IWL<27858> A_IWL<27857> A_IWL<27856> A_IWL<27855> A_IWL<27854> A_IWL<27853> A_IWL<27852> A_IWL<27851> A_IWL<27850> A_IWL<27849> A_IWL<27848> A_IWL<27847> A_IWL<27846> A_IWL<27845> A_IWL<27844> A_IWL<27843> A_IWL<27842> A_IWL<27841> A_IWL<27840> A_IWL<27839> A_IWL<27838> A_IWL<27837> A_IWL<27836> A_IWL<27835> A_IWL<27834> A_IWL<27833> A_IWL<27832> A_IWL<27831> A_IWL<27830> A_IWL<27829> A_IWL<27828> A_IWL<27827> A_IWL<27826> A_IWL<27825> A_IWL<27824> A_IWL<27823> A_IWL<27822> A_IWL<27821> A_IWL<27820> A_IWL<27819> A_IWL<27818> A_IWL<27817> A_IWL<27816> A_IWL<27815> A_IWL<27814> A_IWL<27813> A_IWL<27812> A_IWL<27811> A_IWL<27810> A_IWL<27809> A_IWL<27808> A_IWL<27807> A_IWL<27806> A_IWL<27805> A_IWL<27804> A_IWL<27803> A_IWL<27802> A_IWL<27801> A_IWL<27800> A_IWL<27799> A_IWL<27798> A_IWL<27797> A_IWL<27796> A_IWL<27795> A_IWL<27794> A_IWL<27793> A_IWL<27792> A_IWL<27791> A_IWL<27790> A_IWL<27789> A_IWL<27788> A_IWL<27787> A_IWL<27786> A_IWL<27785> A_IWL<27784> A_IWL<27783> A_IWL<27782> A_IWL<27781> A_IWL<27780> A_IWL<27779> A_IWL<27778> A_IWL<27777> A_IWL<27776> A_IWL<27775> A_IWL<27774> A_IWL<27773> A_IWL<27772> A_IWL<27771> A_IWL<27770> A_IWL<27769> A_IWL<27768> A_IWL<27767> A_IWL<27766> A_IWL<27765> A_IWL<27764> A_IWL<27763> A_IWL<27762> A_IWL<27761> A_IWL<27760> A_IWL<27759> A_IWL<27758> A_IWL<27757> A_IWL<27756> A_IWL<27755> A_IWL<27754> A_IWL<27753> A_IWL<27752> A_IWL<27751> A_IWL<27750> A_IWL<27749> A_IWL<27748> A_IWL<27747> A_IWL<27746> A_IWL<27745> A_IWL<27744> A_IWL<27743> A_IWL<27742> A_IWL<27741> A_IWL<27740> A_IWL<27739> A_IWL<27738> A_IWL<27737> A_IWL<27736> A_IWL<27735> A_IWL<27734> A_IWL<27733> A_IWL<27732> A_IWL<27731> A_IWL<27730> A_IWL<27729> A_IWL<27728> A_IWL<27727> A_IWL<27726> A_IWL<27725> A_IWL<27724> A_IWL<27723> A_IWL<27722> A_IWL<27721> A_IWL<27720> A_IWL<27719> A_IWL<27718> A_IWL<27717> A_IWL<27716> A_IWL<27715> A_IWL<27714> A_IWL<27713> A_IWL<27712> A_IWL<27711> A_IWL<27710> A_IWL<27709> A_IWL<27708> A_IWL<27707> A_IWL<27706> A_IWL<27705> A_IWL<27704> A_IWL<27703> A_IWL<27702> A_IWL<27701> A_IWL<27700> A_IWL<27699> A_IWL<27698> A_IWL<27697> A_IWL<27696> A_IWL<27695> A_IWL<27694> A_IWL<27693> A_IWL<27692> A_IWL<27691> A_IWL<27690> A_IWL<27689> A_IWL<27688> A_IWL<27687> A_IWL<27686> A_IWL<27685> A_IWL<27684> A_IWL<27683> A_IWL<27682> A_IWL<27681> A_IWL<27680> A_IWL<27679> A_IWL<27678> A_IWL<27677> A_IWL<27676> A_IWL<27675> A_IWL<27674> A_IWL<27673> A_IWL<27672> A_IWL<27671> A_IWL<27670> A_IWL<27669> A_IWL<27668> A_IWL<27667> A_IWL<27666> A_IWL<27665> A_IWL<27664> A_IWL<27663> A_IWL<27662> A_IWL<27661> A_IWL<27660> A_IWL<27659> A_IWL<27658> A_IWL<27657> A_IWL<27656> A_IWL<27655> A_IWL<27654> A_IWL<27653> A_IWL<27652> A_IWL<27651> A_IWL<27650> A_IWL<27649> A_IWL<27648> A_IWL<28671> A_IWL<28670> A_IWL<28669> A_IWL<28668> A_IWL<28667> A_IWL<28666> A_IWL<28665> A_IWL<28664> A_IWL<28663> A_IWL<28662> A_IWL<28661> A_IWL<28660> A_IWL<28659> A_IWL<28658> A_IWL<28657> A_IWL<28656> A_IWL<28655> A_IWL<28654> A_IWL<28653> A_IWL<28652> A_IWL<28651> A_IWL<28650> A_IWL<28649> A_IWL<28648> A_IWL<28647> A_IWL<28646> A_IWL<28645> A_IWL<28644> A_IWL<28643> A_IWL<28642> A_IWL<28641> A_IWL<28640> A_IWL<28639> A_IWL<28638> A_IWL<28637> A_IWL<28636> A_IWL<28635> A_IWL<28634> A_IWL<28633> A_IWL<28632> A_IWL<28631> A_IWL<28630> A_IWL<28629> A_IWL<28628> A_IWL<28627> A_IWL<28626> A_IWL<28625> A_IWL<28624> A_IWL<28623> A_IWL<28622> A_IWL<28621> A_IWL<28620> A_IWL<28619> A_IWL<28618> A_IWL<28617> A_IWL<28616> A_IWL<28615> A_IWL<28614> A_IWL<28613> A_IWL<28612> A_IWL<28611> A_IWL<28610> A_IWL<28609> A_IWL<28608> A_IWL<28607> A_IWL<28606> A_IWL<28605> A_IWL<28604> A_IWL<28603> A_IWL<28602> A_IWL<28601> A_IWL<28600> A_IWL<28599> A_IWL<28598> A_IWL<28597> A_IWL<28596> A_IWL<28595> A_IWL<28594> A_IWL<28593> A_IWL<28592> A_IWL<28591> A_IWL<28590> A_IWL<28589> A_IWL<28588> A_IWL<28587> A_IWL<28586> A_IWL<28585> A_IWL<28584> A_IWL<28583> A_IWL<28582> A_IWL<28581> A_IWL<28580> A_IWL<28579> A_IWL<28578> A_IWL<28577> A_IWL<28576> A_IWL<28575> A_IWL<28574> A_IWL<28573> A_IWL<28572> A_IWL<28571> A_IWL<28570> A_IWL<28569> A_IWL<28568> A_IWL<28567> A_IWL<28566> A_IWL<28565> A_IWL<28564> A_IWL<28563> A_IWL<28562> A_IWL<28561> A_IWL<28560> A_IWL<28559> A_IWL<28558> A_IWL<28557> A_IWL<28556> A_IWL<28555> A_IWL<28554> A_IWL<28553> A_IWL<28552> A_IWL<28551> A_IWL<28550> A_IWL<28549> A_IWL<28548> A_IWL<28547> A_IWL<28546> A_IWL<28545> A_IWL<28544> A_IWL<28543> A_IWL<28542> A_IWL<28541> A_IWL<28540> A_IWL<28539> A_IWL<28538> A_IWL<28537> A_IWL<28536> A_IWL<28535> A_IWL<28534> A_IWL<28533> A_IWL<28532> A_IWL<28531> A_IWL<28530> A_IWL<28529> A_IWL<28528> A_IWL<28527> A_IWL<28526> A_IWL<28525> A_IWL<28524> A_IWL<28523> A_IWL<28522> A_IWL<28521> A_IWL<28520> A_IWL<28519> A_IWL<28518> A_IWL<28517> A_IWL<28516> A_IWL<28515> A_IWL<28514> A_IWL<28513> A_IWL<28512> A_IWL<28511> A_IWL<28510> A_IWL<28509> A_IWL<28508> A_IWL<28507> A_IWL<28506> A_IWL<28505> A_IWL<28504> A_IWL<28503> A_IWL<28502> A_IWL<28501> A_IWL<28500> A_IWL<28499> A_IWL<28498> A_IWL<28497> A_IWL<28496> A_IWL<28495> A_IWL<28494> A_IWL<28493> A_IWL<28492> A_IWL<28491> A_IWL<28490> A_IWL<28489> A_IWL<28488> A_IWL<28487> A_IWL<28486> A_IWL<28485> A_IWL<28484> A_IWL<28483> A_IWL<28482> A_IWL<28481> A_IWL<28480> A_IWL<28479> A_IWL<28478> A_IWL<28477> A_IWL<28476> A_IWL<28475> A_IWL<28474> A_IWL<28473> A_IWL<28472> A_IWL<28471> A_IWL<28470> A_IWL<28469> A_IWL<28468> A_IWL<28467> A_IWL<28466> A_IWL<28465> A_IWL<28464> A_IWL<28463> A_IWL<28462> A_IWL<28461> A_IWL<28460> A_IWL<28459> A_IWL<28458> A_IWL<28457> A_IWL<28456> A_IWL<28455> A_IWL<28454> A_IWL<28453> A_IWL<28452> A_IWL<28451> A_IWL<28450> A_IWL<28449> A_IWL<28448> A_IWL<28447> A_IWL<28446> A_IWL<28445> A_IWL<28444> A_IWL<28443> A_IWL<28442> A_IWL<28441> A_IWL<28440> A_IWL<28439> A_IWL<28438> A_IWL<28437> A_IWL<28436> A_IWL<28435> A_IWL<28434> A_IWL<28433> A_IWL<28432> A_IWL<28431> A_IWL<28430> A_IWL<28429> A_IWL<28428> A_IWL<28427> A_IWL<28426> A_IWL<28425> A_IWL<28424> A_IWL<28423> A_IWL<28422> A_IWL<28421> A_IWL<28420> A_IWL<28419> A_IWL<28418> A_IWL<28417> A_IWL<28416> A_IWL<28415> A_IWL<28414> A_IWL<28413> A_IWL<28412> A_IWL<28411> A_IWL<28410> A_IWL<28409> A_IWL<28408> A_IWL<28407> A_IWL<28406> A_IWL<28405> A_IWL<28404> A_IWL<28403> A_IWL<28402> A_IWL<28401> A_IWL<28400> A_IWL<28399> A_IWL<28398> A_IWL<28397> A_IWL<28396> A_IWL<28395> A_IWL<28394> A_IWL<28393> A_IWL<28392> A_IWL<28391> A_IWL<28390> A_IWL<28389> A_IWL<28388> A_IWL<28387> A_IWL<28386> A_IWL<28385> A_IWL<28384> A_IWL<28383> A_IWL<28382> A_IWL<28381> A_IWL<28380> A_IWL<28379> A_IWL<28378> A_IWL<28377> A_IWL<28376> A_IWL<28375> A_IWL<28374> A_IWL<28373> A_IWL<28372> A_IWL<28371> A_IWL<28370> A_IWL<28369> A_IWL<28368> A_IWL<28367> A_IWL<28366> A_IWL<28365> A_IWL<28364> A_IWL<28363> A_IWL<28362> A_IWL<28361> A_IWL<28360> A_IWL<28359> A_IWL<28358> A_IWL<28357> A_IWL<28356> A_IWL<28355> A_IWL<28354> A_IWL<28353> A_IWL<28352> A_IWL<28351> A_IWL<28350> A_IWL<28349> A_IWL<28348> A_IWL<28347> A_IWL<28346> A_IWL<28345> A_IWL<28344> A_IWL<28343> A_IWL<28342> A_IWL<28341> A_IWL<28340> A_IWL<28339> A_IWL<28338> A_IWL<28337> A_IWL<28336> A_IWL<28335> A_IWL<28334> A_IWL<28333> A_IWL<28332> A_IWL<28331> A_IWL<28330> A_IWL<28329> A_IWL<28328> A_IWL<28327> A_IWL<28326> A_IWL<28325> A_IWL<28324> A_IWL<28323> A_IWL<28322> A_IWL<28321> A_IWL<28320> A_IWL<28319> A_IWL<28318> A_IWL<28317> A_IWL<28316> A_IWL<28315> A_IWL<28314> A_IWL<28313> A_IWL<28312> A_IWL<28311> A_IWL<28310> A_IWL<28309> A_IWL<28308> A_IWL<28307> A_IWL<28306> A_IWL<28305> A_IWL<28304> A_IWL<28303> A_IWL<28302> A_IWL<28301> A_IWL<28300> A_IWL<28299> A_IWL<28298> A_IWL<28297> A_IWL<28296> A_IWL<28295> A_IWL<28294> A_IWL<28293> A_IWL<28292> A_IWL<28291> A_IWL<28290> A_IWL<28289> A_IWL<28288> A_IWL<28287> A_IWL<28286> A_IWL<28285> A_IWL<28284> A_IWL<28283> A_IWL<28282> A_IWL<28281> A_IWL<28280> A_IWL<28279> A_IWL<28278> A_IWL<28277> A_IWL<28276> A_IWL<28275> A_IWL<28274> A_IWL<28273> A_IWL<28272> A_IWL<28271> A_IWL<28270> A_IWL<28269> A_IWL<28268> A_IWL<28267> A_IWL<28266> A_IWL<28265> A_IWL<28264> A_IWL<28263> A_IWL<28262> A_IWL<28261> A_IWL<28260> A_IWL<28259> A_IWL<28258> A_IWL<28257> A_IWL<28256> A_IWL<28255> A_IWL<28254> A_IWL<28253> A_IWL<28252> A_IWL<28251> A_IWL<28250> A_IWL<28249> A_IWL<28248> A_IWL<28247> A_IWL<28246> A_IWL<28245> A_IWL<28244> A_IWL<28243> A_IWL<28242> A_IWL<28241> A_IWL<28240> A_IWL<28239> A_IWL<28238> A_IWL<28237> A_IWL<28236> A_IWL<28235> A_IWL<28234> A_IWL<28233> A_IWL<28232> A_IWL<28231> A_IWL<28230> A_IWL<28229> A_IWL<28228> A_IWL<28227> A_IWL<28226> A_IWL<28225> A_IWL<28224> A_IWL<28223> A_IWL<28222> A_IWL<28221> A_IWL<28220> A_IWL<28219> A_IWL<28218> A_IWL<28217> A_IWL<28216> A_IWL<28215> A_IWL<28214> A_IWL<28213> A_IWL<28212> A_IWL<28211> A_IWL<28210> A_IWL<28209> A_IWL<28208> A_IWL<28207> A_IWL<28206> A_IWL<28205> A_IWL<28204> A_IWL<28203> A_IWL<28202> A_IWL<28201> A_IWL<28200> A_IWL<28199> A_IWL<28198> A_IWL<28197> A_IWL<28196> A_IWL<28195> A_IWL<28194> A_IWL<28193> A_IWL<28192> A_IWL<28191> A_IWL<28190> A_IWL<28189> A_IWL<28188> A_IWL<28187> A_IWL<28186> A_IWL<28185> A_IWL<28184> A_IWL<28183> A_IWL<28182> A_IWL<28181> A_IWL<28180> A_IWL<28179> A_IWL<28178> A_IWL<28177> A_IWL<28176> A_IWL<28175> A_IWL<28174> A_IWL<28173> A_IWL<28172> A_IWL<28171> A_IWL<28170> A_IWL<28169> A_IWL<28168> A_IWL<28167> A_IWL<28166> A_IWL<28165> A_IWL<28164> A_IWL<28163> A_IWL<28162> A_IWL<28161> A_IWL<28160> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<54> A_BLC<109> A_BLC<108> A_BLC_TOP<109> A_BLC_TOP<108> A_BLT<109> A_BLT<108> A_BLT_TOP<109> A_BLT_TOP<108> A_IWL<27647> A_IWL<27646> A_IWL<27645> A_IWL<27644> A_IWL<27643> A_IWL<27642> A_IWL<27641> A_IWL<27640> A_IWL<27639> A_IWL<27638> A_IWL<27637> A_IWL<27636> A_IWL<27635> A_IWL<27634> A_IWL<27633> A_IWL<27632> A_IWL<27631> A_IWL<27630> A_IWL<27629> A_IWL<27628> A_IWL<27627> A_IWL<27626> A_IWL<27625> A_IWL<27624> A_IWL<27623> A_IWL<27622> A_IWL<27621> A_IWL<27620> A_IWL<27619> A_IWL<27618> A_IWL<27617> A_IWL<27616> A_IWL<27615> A_IWL<27614> A_IWL<27613> A_IWL<27612> A_IWL<27611> A_IWL<27610> A_IWL<27609> A_IWL<27608> A_IWL<27607> A_IWL<27606> A_IWL<27605> A_IWL<27604> A_IWL<27603> A_IWL<27602> A_IWL<27601> A_IWL<27600> A_IWL<27599> A_IWL<27598> A_IWL<27597> A_IWL<27596> A_IWL<27595> A_IWL<27594> A_IWL<27593> A_IWL<27592> A_IWL<27591> A_IWL<27590> A_IWL<27589> A_IWL<27588> A_IWL<27587> A_IWL<27586> A_IWL<27585> A_IWL<27584> A_IWL<27583> A_IWL<27582> A_IWL<27581> A_IWL<27580> A_IWL<27579> A_IWL<27578> A_IWL<27577> A_IWL<27576> A_IWL<27575> A_IWL<27574> A_IWL<27573> A_IWL<27572> A_IWL<27571> A_IWL<27570> A_IWL<27569> A_IWL<27568> A_IWL<27567> A_IWL<27566> A_IWL<27565> A_IWL<27564> A_IWL<27563> A_IWL<27562> A_IWL<27561> A_IWL<27560> A_IWL<27559> A_IWL<27558> A_IWL<27557> A_IWL<27556> A_IWL<27555> A_IWL<27554> A_IWL<27553> A_IWL<27552> A_IWL<27551> A_IWL<27550> A_IWL<27549> A_IWL<27548> A_IWL<27547> A_IWL<27546> A_IWL<27545> A_IWL<27544> A_IWL<27543> A_IWL<27542> A_IWL<27541> A_IWL<27540> A_IWL<27539> A_IWL<27538> A_IWL<27537> A_IWL<27536> A_IWL<27535> A_IWL<27534> A_IWL<27533> A_IWL<27532> A_IWL<27531> A_IWL<27530> A_IWL<27529> A_IWL<27528> A_IWL<27527> A_IWL<27526> A_IWL<27525> A_IWL<27524> A_IWL<27523> A_IWL<27522> A_IWL<27521> A_IWL<27520> A_IWL<27519> A_IWL<27518> A_IWL<27517> A_IWL<27516> A_IWL<27515> A_IWL<27514> A_IWL<27513> A_IWL<27512> A_IWL<27511> A_IWL<27510> A_IWL<27509> A_IWL<27508> A_IWL<27507> A_IWL<27506> A_IWL<27505> A_IWL<27504> A_IWL<27503> A_IWL<27502> A_IWL<27501> A_IWL<27500> A_IWL<27499> A_IWL<27498> A_IWL<27497> A_IWL<27496> A_IWL<27495> A_IWL<27494> A_IWL<27493> A_IWL<27492> A_IWL<27491> A_IWL<27490> A_IWL<27489> A_IWL<27488> A_IWL<27487> A_IWL<27486> A_IWL<27485> A_IWL<27484> A_IWL<27483> A_IWL<27482> A_IWL<27481> A_IWL<27480> A_IWL<27479> A_IWL<27478> A_IWL<27477> A_IWL<27476> A_IWL<27475> A_IWL<27474> A_IWL<27473> A_IWL<27472> A_IWL<27471> A_IWL<27470> A_IWL<27469> A_IWL<27468> A_IWL<27467> A_IWL<27466> A_IWL<27465> A_IWL<27464> A_IWL<27463> A_IWL<27462> A_IWL<27461> A_IWL<27460> A_IWL<27459> A_IWL<27458> A_IWL<27457> A_IWL<27456> A_IWL<27455> A_IWL<27454> A_IWL<27453> A_IWL<27452> A_IWL<27451> A_IWL<27450> A_IWL<27449> A_IWL<27448> A_IWL<27447> A_IWL<27446> A_IWL<27445> A_IWL<27444> A_IWL<27443> A_IWL<27442> A_IWL<27441> A_IWL<27440> A_IWL<27439> A_IWL<27438> A_IWL<27437> A_IWL<27436> A_IWL<27435> A_IWL<27434> A_IWL<27433> A_IWL<27432> A_IWL<27431> A_IWL<27430> A_IWL<27429> A_IWL<27428> A_IWL<27427> A_IWL<27426> A_IWL<27425> A_IWL<27424> A_IWL<27423> A_IWL<27422> A_IWL<27421> A_IWL<27420> A_IWL<27419> A_IWL<27418> A_IWL<27417> A_IWL<27416> A_IWL<27415> A_IWL<27414> A_IWL<27413> A_IWL<27412> A_IWL<27411> A_IWL<27410> A_IWL<27409> A_IWL<27408> A_IWL<27407> A_IWL<27406> A_IWL<27405> A_IWL<27404> A_IWL<27403> A_IWL<27402> A_IWL<27401> A_IWL<27400> A_IWL<27399> A_IWL<27398> A_IWL<27397> A_IWL<27396> A_IWL<27395> A_IWL<27394> A_IWL<27393> A_IWL<27392> A_IWL<27391> A_IWL<27390> A_IWL<27389> A_IWL<27388> A_IWL<27387> A_IWL<27386> A_IWL<27385> A_IWL<27384> A_IWL<27383> A_IWL<27382> A_IWL<27381> A_IWL<27380> A_IWL<27379> A_IWL<27378> A_IWL<27377> A_IWL<27376> A_IWL<27375> A_IWL<27374> A_IWL<27373> A_IWL<27372> A_IWL<27371> A_IWL<27370> A_IWL<27369> A_IWL<27368> A_IWL<27367> A_IWL<27366> A_IWL<27365> A_IWL<27364> A_IWL<27363> A_IWL<27362> A_IWL<27361> A_IWL<27360> A_IWL<27359> A_IWL<27358> A_IWL<27357> A_IWL<27356> A_IWL<27355> A_IWL<27354> A_IWL<27353> A_IWL<27352> A_IWL<27351> A_IWL<27350> A_IWL<27349> A_IWL<27348> A_IWL<27347> A_IWL<27346> A_IWL<27345> A_IWL<27344> A_IWL<27343> A_IWL<27342> A_IWL<27341> A_IWL<27340> A_IWL<27339> A_IWL<27338> A_IWL<27337> A_IWL<27336> A_IWL<27335> A_IWL<27334> A_IWL<27333> A_IWL<27332> A_IWL<27331> A_IWL<27330> A_IWL<27329> A_IWL<27328> A_IWL<27327> A_IWL<27326> A_IWL<27325> A_IWL<27324> A_IWL<27323> A_IWL<27322> A_IWL<27321> A_IWL<27320> A_IWL<27319> A_IWL<27318> A_IWL<27317> A_IWL<27316> A_IWL<27315> A_IWL<27314> A_IWL<27313> A_IWL<27312> A_IWL<27311> A_IWL<27310> A_IWL<27309> A_IWL<27308> A_IWL<27307> A_IWL<27306> A_IWL<27305> A_IWL<27304> A_IWL<27303> A_IWL<27302> A_IWL<27301> A_IWL<27300> A_IWL<27299> A_IWL<27298> A_IWL<27297> A_IWL<27296> A_IWL<27295> A_IWL<27294> A_IWL<27293> A_IWL<27292> A_IWL<27291> A_IWL<27290> A_IWL<27289> A_IWL<27288> A_IWL<27287> A_IWL<27286> A_IWL<27285> A_IWL<27284> A_IWL<27283> A_IWL<27282> A_IWL<27281> A_IWL<27280> A_IWL<27279> A_IWL<27278> A_IWL<27277> A_IWL<27276> A_IWL<27275> A_IWL<27274> A_IWL<27273> A_IWL<27272> A_IWL<27271> A_IWL<27270> A_IWL<27269> A_IWL<27268> A_IWL<27267> A_IWL<27266> A_IWL<27265> A_IWL<27264> A_IWL<27263> A_IWL<27262> A_IWL<27261> A_IWL<27260> A_IWL<27259> A_IWL<27258> A_IWL<27257> A_IWL<27256> A_IWL<27255> A_IWL<27254> A_IWL<27253> A_IWL<27252> A_IWL<27251> A_IWL<27250> A_IWL<27249> A_IWL<27248> A_IWL<27247> A_IWL<27246> A_IWL<27245> A_IWL<27244> A_IWL<27243> A_IWL<27242> A_IWL<27241> A_IWL<27240> A_IWL<27239> A_IWL<27238> A_IWL<27237> A_IWL<27236> A_IWL<27235> A_IWL<27234> A_IWL<27233> A_IWL<27232> A_IWL<27231> A_IWL<27230> A_IWL<27229> A_IWL<27228> A_IWL<27227> A_IWL<27226> A_IWL<27225> A_IWL<27224> A_IWL<27223> A_IWL<27222> A_IWL<27221> A_IWL<27220> A_IWL<27219> A_IWL<27218> A_IWL<27217> A_IWL<27216> A_IWL<27215> A_IWL<27214> A_IWL<27213> A_IWL<27212> A_IWL<27211> A_IWL<27210> A_IWL<27209> A_IWL<27208> A_IWL<27207> A_IWL<27206> A_IWL<27205> A_IWL<27204> A_IWL<27203> A_IWL<27202> A_IWL<27201> A_IWL<27200> A_IWL<27199> A_IWL<27198> A_IWL<27197> A_IWL<27196> A_IWL<27195> A_IWL<27194> A_IWL<27193> A_IWL<27192> A_IWL<27191> A_IWL<27190> A_IWL<27189> A_IWL<27188> A_IWL<27187> A_IWL<27186> A_IWL<27185> A_IWL<27184> A_IWL<27183> A_IWL<27182> A_IWL<27181> A_IWL<27180> A_IWL<27179> A_IWL<27178> A_IWL<27177> A_IWL<27176> A_IWL<27175> A_IWL<27174> A_IWL<27173> A_IWL<27172> A_IWL<27171> A_IWL<27170> A_IWL<27169> A_IWL<27168> A_IWL<27167> A_IWL<27166> A_IWL<27165> A_IWL<27164> A_IWL<27163> A_IWL<27162> A_IWL<27161> A_IWL<27160> A_IWL<27159> A_IWL<27158> A_IWL<27157> A_IWL<27156> A_IWL<27155> A_IWL<27154> A_IWL<27153> A_IWL<27152> A_IWL<27151> A_IWL<27150> A_IWL<27149> A_IWL<27148> A_IWL<27147> A_IWL<27146> A_IWL<27145> A_IWL<27144> A_IWL<27143> A_IWL<27142> A_IWL<27141> A_IWL<27140> A_IWL<27139> A_IWL<27138> A_IWL<27137> A_IWL<27136> A_IWL<28159> A_IWL<28158> A_IWL<28157> A_IWL<28156> A_IWL<28155> A_IWL<28154> A_IWL<28153> A_IWL<28152> A_IWL<28151> A_IWL<28150> A_IWL<28149> A_IWL<28148> A_IWL<28147> A_IWL<28146> A_IWL<28145> A_IWL<28144> A_IWL<28143> A_IWL<28142> A_IWL<28141> A_IWL<28140> A_IWL<28139> A_IWL<28138> A_IWL<28137> A_IWL<28136> A_IWL<28135> A_IWL<28134> A_IWL<28133> A_IWL<28132> A_IWL<28131> A_IWL<28130> A_IWL<28129> A_IWL<28128> A_IWL<28127> A_IWL<28126> A_IWL<28125> A_IWL<28124> A_IWL<28123> A_IWL<28122> A_IWL<28121> A_IWL<28120> A_IWL<28119> A_IWL<28118> A_IWL<28117> A_IWL<28116> A_IWL<28115> A_IWL<28114> A_IWL<28113> A_IWL<28112> A_IWL<28111> A_IWL<28110> A_IWL<28109> A_IWL<28108> A_IWL<28107> A_IWL<28106> A_IWL<28105> A_IWL<28104> A_IWL<28103> A_IWL<28102> A_IWL<28101> A_IWL<28100> A_IWL<28099> A_IWL<28098> A_IWL<28097> A_IWL<28096> A_IWL<28095> A_IWL<28094> A_IWL<28093> A_IWL<28092> A_IWL<28091> A_IWL<28090> A_IWL<28089> A_IWL<28088> A_IWL<28087> A_IWL<28086> A_IWL<28085> A_IWL<28084> A_IWL<28083> A_IWL<28082> A_IWL<28081> A_IWL<28080> A_IWL<28079> A_IWL<28078> A_IWL<28077> A_IWL<28076> A_IWL<28075> A_IWL<28074> A_IWL<28073> A_IWL<28072> A_IWL<28071> A_IWL<28070> A_IWL<28069> A_IWL<28068> A_IWL<28067> A_IWL<28066> A_IWL<28065> A_IWL<28064> A_IWL<28063> A_IWL<28062> A_IWL<28061> A_IWL<28060> A_IWL<28059> A_IWL<28058> A_IWL<28057> A_IWL<28056> A_IWL<28055> A_IWL<28054> A_IWL<28053> A_IWL<28052> A_IWL<28051> A_IWL<28050> A_IWL<28049> A_IWL<28048> A_IWL<28047> A_IWL<28046> A_IWL<28045> A_IWL<28044> A_IWL<28043> A_IWL<28042> A_IWL<28041> A_IWL<28040> A_IWL<28039> A_IWL<28038> A_IWL<28037> A_IWL<28036> A_IWL<28035> A_IWL<28034> A_IWL<28033> A_IWL<28032> A_IWL<28031> A_IWL<28030> A_IWL<28029> A_IWL<28028> A_IWL<28027> A_IWL<28026> A_IWL<28025> A_IWL<28024> A_IWL<28023> A_IWL<28022> A_IWL<28021> A_IWL<28020> A_IWL<28019> A_IWL<28018> A_IWL<28017> A_IWL<28016> A_IWL<28015> A_IWL<28014> A_IWL<28013> A_IWL<28012> A_IWL<28011> A_IWL<28010> A_IWL<28009> A_IWL<28008> A_IWL<28007> A_IWL<28006> A_IWL<28005> A_IWL<28004> A_IWL<28003> A_IWL<28002> A_IWL<28001> A_IWL<28000> A_IWL<27999> A_IWL<27998> A_IWL<27997> A_IWL<27996> A_IWL<27995> A_IWL<27994> A_IWL<27993> A_IWL<27992> A_IWL<27991> A_IWL<27990> A_IWL<27989> A_IWL<27988> A_IWL<27987> A_IWL<27986> A_IWL<27985> A_IWL<27984> A_IWL<27983> A_IWL<27982> A_IWL<27981> A_IWL<27980> A_IWL<27979> A_IWL<27978> A_IWL<27977> A_IWL<27976> A_IWL<27975> A_IWL<27974> A_IWL<27973> A_IWL<27972> A_IWL<27971> A_IWL<27970> A_IWL<27969> A_IWL<27968> A_IWL<27967> A_IWL<27966> A_IWL<27965> A_IWL<27964> A_IWL<27963> A_IWL<27962> A_IWL<27961> A_IWL<27960> A_IWL<27959> A_IWL<27958> A_IWL<27957> A_IWL<27956> A_IWL<27955> A_IWL<27954> A_IWL<27953> A_IWL<27952> A_IWL<27951> A_IWL<27950> A_IWL<27949> A_IWL<27948> A_IWL<27947> A_IWL<27946> A_IWL<27945> A_IWL<27944> A_IWL<27943> A_IWL<27942> A_IWL<27941> A_IWL<27940> A_IWL<27939> A_IWL<27938> A_IWL<27937> A_IWL<27936> A_IWL<27935> A_IWL<27934> A_IWL<27933> A_IWL<27932> A_IWL<27931> A_IWL<27930> A_IWL<27929> A_IWL<27928> A_IWL<27927> A_IWL<27926> A_IWL<27925> A_IWL<27924> A_IWL<27923> A_IWL<27922> A_IWL<27921> A_IWL<27920> A_IWL<27919> A_IWL<27918> A_IWL<27917> A_IWL<27916> A_IWL<27915> A_IWL<27914> A_IWL<27913> A_IWL<27912> A_IWL<27911> A_IWL<27910> A_IWL<27909> A_IWL<27908> A_IWL<27907> A_IWL<27906> A_IWL<27905> A_IWL<27904> A_IWL<27903> A_IWL<27902> A_IWL<27901> A_IWL<27900> A_IWL<27899> A_IWL<27898> A_IWL<27897> A_IWL<27896> A_IWL<27895> A_IWL<27894> A_IWL<27893> A_IWL<27892> A_IWL<27891> A_IWL<27890> A_IWL<27889> A_IWL<27888> A_IWL<27887> A_IWL<27886> A_IWL<27885> A_IWL<27884> A_IWL<27883> A_IWL<27882> A_IWL<27881> A_IWL<27880> A_IWL<27879> A_IWL<27878> A_IWL<27877> A_IWL<27876> A_IWL<27875> A_IWL<27874> A_IWL<27873> A_IWL<27872> A_IWL<27871> A_IWL<27870> A_IWL<27869> A_IWL<27868> A_IWL<27867> A_IWL<27866> A_IWL<27865> A_IWL<27864> A_IWL<27863> A_IWL<27862> A_IWL<27861> A_IWL<27860> A_IWL<27859> A_IWL<27858> A_IWL<27857> A_IWL<27856> A_IWL<27855> A_IWL<27854> A_IWL<27853> A_IWL<27852> A_IWL<27851> A_IWL<27850> A_IWL<27849> A_IWL<27848> A_IWL<27847> A_IWL<27846> A_IWL<27845> A_IWL<27844> A_IWL<27843> A_IWL<27842> A_IWL<27841> A_IWL<27840> A_IWL<27839> A_IWL<27838> A_IWL<27837> A_IWL<27836> A_IWL<27835> A_IWL<27834> A_IWL<27833> A_IWL<27832> A_IWL<27831> A_IWL<27830> A_IWL<27829> A_IWL<27828> A_IWL<27827> A_IWL<27826> A_IWL<27825> A_IWL<27824> A_IWL<27823> A_IWL<27822> A_IWL<27821> A_IWL<27820> A_IWL<27819> A_IWL<27818> A_IWL<27817> A_IWL<27816> A_IWL<27815> A_IWL<27814> A_IWL<27813> A_IWL<27812> A_IWL<27811> A_IWL<27810> A_IWL<27809> A_IWL<27808> A_IWL<27807> A_IWL<27806> A_IWL<27805> A_IWL<27804> A_IWL<27803> A_IWL<27802> A_IWL<27801> A_IWL<27800> A_IWL<27799> A_IWL<27798> A_IWL<27797> A_IWL<27796> A_IWL<27795> A_IWL<27794> A_IWL<27793> A_IWL<27792> A_IWL<27791> A_IWL<27790> A_IWL<27789> A_IWL<27788> A_IWL<27787> A_IWL<27786> A_IWL<27785> A_IWL<27784> A_IWL<27783> A_IWL<27782> A_IWL<27781> A_IWL<27780> A_IWL<27779> A_IWL<27778> A_IWL<27777> A_IWL<27776> A_IWL<27775> A_IWL<27774> A_IWL<27773> A_IWL<27772> A_IWL<27771> A_IWL<27770> A_IWL<27769> A_IWL<27768> A_IWL<27767> A_IWL<27766> A_IWL<27765> A_IWL<27764> A_IWL<27763> A_IWL<27762> A_IWL<27761> A_IWL<27760> A_IWL<27759> A_IWL<27758> A_IWL<27757> A_IWL<27756> A_IWL<27755> A_IWL<27754> A_IWL<27753> A_IWL<27752> A_IWL<27751> A_IWL<27750> A_IWL<27749> A_IWL<27748> A_IWL<27747> A_IWL<27746> A_IWL<27745> A_IWL<27744> A_IWL<27743> A_IWL<27742> A_IWL<27741> A_IWL<27740> A_IWL<27739> A_IWL<27738> A_IWL<27737> A_IWL<27736> A_IWL<27735> A_IWL<27734> A_IWL<27733> A_IWL<27732> A_IWL<27731> A_IWL<27730> A_IWL<27729> A_IWL<27728> A_IWL<27727> A_IWL<27726> A_IWL<27725> A_IWL<27724> A_IWL<27723> A_IWL<27722> A_IWL<27721> A_IWL<27720> A_IWL<27719> A_IWL<27718> A_IWL<27717> A_IWL<27716> A_IWL<27715> A_IWL<27714> A_IWL<27713> A_IWL<27712> A_IWL<27711> A_IWL<27710> A_IWL<27709> A_IWL<27708> A_IWL<27707> A_IWL<27706> A_IWL<27705> A_IWL<27704> A_IWL<27703> A_IWL<27702> A_IWL<27701> A_IWL<27700> A_IWL<27699> A_IWL<27698> A_IWL<27697> A_IWL<27696> A_IWL<27695> A_IWL<27694> A_IWL<27693> A_IWL<27692> A_IWL<27691> A_IWL<27690> A_IWL<27689> A_IWL<27688> A_IWL<27687> A_IWL<27686> A_IWL<27685> A_IWL<27684> A_IWL<27683> A_IWL<27682> A_IWL<27681> A_IWL<27680> A_IWL<27679> A_IWL<27678> A_IWL<27677> A_IWL<27676> A_IWL<27675> A_IWL<27674> A_IWL<27673> A_IWL<27672> A_IWL<27671> A_IWL<27670> A_IWL<27669> A_IWL<27668> A_IWL<27667> A_IWL<27666> A_IWL<27665> A_IWL<27664> A_IWL<27663> A_IWL<27662> A_IWL<27661> A_IWL<27660> A_IWL<27659> A_IWL<27658> A_IWL<27657> A_IWL<27656> A_IWL<27655> A_IWL<27654> A_IWL<27653> A_IWL<27652> A_IWL<27651> A_IWL<27650> A_IWL<27649> A_IWL<27648> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<53> A_BLC<107> A_BLC<106> A_BLC_TOP<107> A_BLC_TOP<106> A_BLT<107> A_BLT<106> A_BLT_TOP<107> A_BLT_TOP<106> A_IWL<27135> A_IWL<27134> A_IWL<27133> A_IWL<27132> A_IWL<27131> A_IWL<27130> A_IWL<27129> A_IWL<27128> A_IWL<27127> A_IWL<27126> A_IWL<27125> A_IWL<27124> A_IWL<27123> A_IWL<27122> A_IWL<27121> A_IWL<27120> A_IWL<27119> A_IWL<27118> A_IWL<27117> A_IWL<27116> A_IWL<27115> A_IWL<27114> A_IWL<27113> A_IWL<27112> A_IWL<27111> A_IWL<27110> A_IWL<27109> A_IWL<27108> A_IWL<27107> A_IWL<27106> A_IWL<27105> A_IWL<27104> A_IWL<27103> A_IWL<27102> A_IWL<27101> A_IWL<27100> A_IWL<27099> A_IWL<27098> A_IWL<27097> A_IWL<27096> A_IWL<27095> A_IWL<27094> A_IWL<27093> A_IWL<27092> A_IWL<27091> A_IWL<27090> A_IWL<27089> A_IWL<27088> A_IWL<27087> A_IWL<27086> A_IWL<27085> A_IWL<27084> A_IWL<27083> A_IWL<27082> A_IWL<27081> A_IWL<27080> A_IWL<27079> A_IWL<27078> A_IWL<27077> A_IWL<27076> A_IWL<27075> A_IWL<27074> A_IWL<27073> A_IWL<27072> A_IWL<27071> A_IWL<27070> A_IWL<27069> A_IWL<27068> A_IWL<27067> A_IWL<27066> A_IWL<27065> A_IWL<27064> A_IWL<27063> A_IWL<27062> A_IWL<27061> A_IWL<27060> A_IWL<27059> A_IWL<27058> A_IWL<27057> A_IWL<27056> A_IWL<27055> A_IWL<27054> A_IWL<27053> A_IWL<27052> A_IWL<27051> A_IWL<27050> A_IWL<27049> A_IWL<27048> A_IWL<27047> A_IWL<27046> A_IWL<27045> A_IWL<27044> A_IWL<27043> A_IWL<27042> A_IWL<27041> A_IWL<27040> A_IWL<27039> A_IWL<27038> A_IWL<27037> A_IWL<27036> A_IWL<27035> A_IWL<27034> A_IWL<27033> A_IWL<27032> A_IWL<27031> A_IWL<27030> A_IWL<27029> A_IWL<27028> A_IWL<27027> A_IWL<27026> A_IWL<27025> A_IWL<27024> A_IWL<27023> A_IWL<27022> A_IWL<27021> A_IWL<27020> A_IWL<27019> A_IWL<27018> A_IWL<27017> A_IWL<27016> A_IWL<27015> A_IWL<27014> A_IWL<27013> A_IWL<27012> A_IWL<27011> A_IWL<27010> A_IWL<27009> A_IWL<27008> A_IWL<27007> A_IWL<27006> A_IWL<27005> A_IWL<27004> A_IWL<27003> A_IWL<27002> A_IWL<27001> A_IWL<27000> A_IWL<26999> A_IWL<26998> A_IWL<26997> A_IWL<26996> A_IWL<26995> A_IWL<26994> A_IWL<26993> A_IWL<26992> A_IWL<26991> A_IWL<26990> A_IWL<26989> A_IWL<26988> A_IWL<26987> A_IWL<26986> A_IWL<26985> A_IWL<26984> A_IWL<26983> A_IWL<26982> A_IWL<26981> A_IWL<26980> A_IWL<26979> A_IWL<26978> A_IWL<26977> A_IWL<26976> A_IWL<26975> A_IWL<26974> A_IWL<26973> A_IWL<26972> A_IWL<26971> A_IWL<26970> A_IWL<26969> A_IWL<26968> A_IWL<26967> A_IWL<26966> A_IWL<26965> A_IWL<26964> A_IWL<26963> A_IWL<26962> A_IWL<26961> A_IWL<26960> A_IWL<26959> A_IWL<26958> A_IWL<26957> A_IWL<26956> A_IWL<26955> A_IWL<26954> A_IWL<26953> A_IWL<26952> A_IWL<26951> A_IWL<26950> A_IWL<26949> A_IWL<26948> A_IWL<26947> A_IWL<26946> A_IWL<26945> A_IWL<26944> A_IWL<26943> A_IWL<26942> A_IWL<26941> A_IWL<26940> A_IWL<26939> A_IWL<26938> A_IWL<26937> A_IWL<26936> A_IWL<26935> A_IWL<26934> A_IWL<26933> A_IWL<26932> A_IWL<26931> A_IWL<26930> A_IWL<26929> A_IWL<26928> A_IWL<26927> A_IWL<26926> A_IWL<26925> A_IWL<26924> A_IWL<26923> A_IWL<26922> A_IWL<26921> A_IWL<26920> A_IWL<26919> A_IWL<26918> A_IWL<26917> A_IWL<26916> A_IWL<26915> A_IWL<26914> A_IWL<26913> A_IWL<26912> A_IWL<26911> A_IWL<26910> A_IWL<26909> A_IWL<26908> A_IWL<26907> A_IWL<26906> A_IWL<26905> A_IWL<26904> A_IWL<26903> A_IWL<26902> A_IWL<26901> A_IWL<26900> A_IWL<26899> A_IWL<26898> A_IWL<26897> A_IWL<26896> A_IWL<26895> A_IWL<26894> A_IWL<26893> A_IWL<26892> A_IWL<26891> A_IWL<26890> A_IWL<26889> A_IWL<26888> A_IWL<26887> A_IWL<26886> A_IWL<26885> A_IWL<26884> A_IWL<26883> A_IWL<26882> A_IWL<26881> A_IWL<26880> A_IWL<26879> A_IWL<26878> A_IWL<26877> A_IWL<26876> A_IWL<26875> A_IWL<26874> A_IWL<26873> A_IWL<26872> A_IWL<26871> A_IWL<26870> A_IWL<26869> A_IWL<26868> A_IWL<26867> A_IWL<26866> A_IWL<26865> A_IWL<26864> A_IWL<26863> A_IWL<26862> A_IWL<26861> A_IWL<26860> A_IWL<26859> A_IWL<26858> A_IWL<26857> A_IWL<26856> A_IWL<26855> A_IWL<26854> A_IWL<26853> A_IWL<26852> A_IWL<26851> A_IWL<26850> A_IWL<26849> A_IWL<26848> A_IWL<26847> A_IWL<26846> A_IWL<26845> A_IWL<26844> A_IWL<26843> A_IWL<26842> A_IWL<26841> A_IWL<26840> A_IWL<26839> A_IWL<26838> A_IWL<26837> A_IWL<26836> A_IWL<26835> A_IWL<26834> A_IWL<26833> A_IWL<26832> A_IWL<26831> A_IWL<26830> A_IWL<26829> A_IWL<26828> A_IWL<26827> A_IWL<26826> A_IWL<26825> A_IWL<26824> A_IWL<26823> A_IWL<26822> A_IWL<26821> A_IWL<26820> A_IWL<26819> A_IWL<26818> A_IWL<26817> A_IWL<26816> A_IWL<26815> A_IWL<26814> A_IWL<26813> A_IWL<26812> A_IWL<26811> A_IWL<26810> A_IWL<26809> A_IWL<26808> A_IWL<26807> A_IWL<26806> A_IWL<26805> A_IWL<26804> A_IWL<26803> A_IWL<26802> A_IWL<26801> A_IWL<26800> A_IWL<26799> A_IWL<26798> A_IWL<26797> A_IWL<26796> A_IWL<26795> A_IWL<26794> A_IWL<26793> A_IWL<26792> A_IWL<26791> A_IWL<26790> A_IWL<26789> A_IWL<26788> A_IWL<26787> A_IWL<26786> A_IWL<26785> A_IWL<26784> A_IWL<26783> A_IWL<26782> A_IWL<26781> A_IWL<26780> A_IWL<26779> A_IWL<26778> A_IWL<26777> A_IWL<26776> A_IWL<26775> A_IWL<26774> A_IWL<26773> A_IWL<26772> A_IWL<26771> A_IWL<26770> A_IWL<26769> A_IWL<26768> A_IWL<26767> A_IWL<26766> A_IWL<26765> A_IWL<26764> A_IWL<26763> A_IWL<26762> A_IWL<26761> A_IWL<26760> A_IWL<26759> A_IWL<26758> A_IWL<26757> A_IWL<26756> A_IWL<26755> A_IWL<26754> A_IWL<26753> A_IWL<26752> A_IWL<26751> A_IWL<26750> A_IWL<26749> A_IWL<26748> A_IWL<26747> A_IWL<26746> A_IWL<26745> A_IWL<26744> A_IWL<26743> A_IWL<26742> A_IWL<26741> A_IWL<26740> A_IWL<26739> A_IWL<26738> A_IWL<26737> A_IWL<26736> A_IWL<26735> A_IWL<26734> A_IWL<26733> A_IWL<26732> A_IWL<26731> A_IWL<26730> A_IWL<26729> A_IWL<26728> A_IWL<26727> A_IWL<26726> A_IWL<26725> A_IWL<26724> A_IWL<26723> A_IWL<26722> A_IWL<26721> A_IWL<26720> A_IWL<26719> A_IWL<26718> A_IWL<26717> A_IWL<26716> A_IWL<26715> A_IWL<26714> A_IWL<26713> A_IWL<26712> A_IWL<26711> A_IWL<26710> A_IWL<26709> A_IWL<26708> A_IWL<26707> A_IWL<26706> A_IWL<26705> A_IWL<26704> A_IWL<26703> A_IWL<26702> A_IWL<26701> A_IWL<26700> A_IWL<26699> A_IWL<26698> A_IWL<26697> A_IWL<26696> A_IWL<26695> A_IWL<26694> A_IWL<26693> A_IWL<26692> A_IWL<26691> A_IWL<26690> A_IWL<26689> A_IWL<26688> A_IWL<26687> A_IWL<26686> A_IWL<26685> A_IWL<26684> A_IWL<26683> A_IWL<26682> A_IWL<26681> A_IWL<26680> A_IWL<26679> A_IWL<26678> A_IWL<26677> A_IWL<26676> A_IWL<26675> A_IWL<26674> A_IWL<26673> A_IWL<26672> A_IWL<26671> A_IWL<26670> A_IWL<26669> A_IWL<26668> A_IWL<26667> A_IWL<26666> A_IWL<26665> A_IWL<26664> A_IWL<26663> A_IWL<26662> A_IWL<26661> A_IWL<26660> A_IWL<26659> A_IWL<26658> A_IWL<26657> A_IWL<26656> A_IWL<26655> A_IWL<26654> A_IWL<26653> A_IWL<26652> A_IWL<26651> A_IWL<26650> A_IWL<26649> A_IWL<26648> A_IWL<26647> A_IWL<26646> A_IWL<26645> A_IWL<26644> A_IWL<26643> A_IWL<26642> A_IWL<26641> A_IWL<26640> A_IWL<26639> A_IWL<26638> A_IWL<26637> A_IWL<26636> A_IWL<26635> A_IWL<26634> A_IWL<26633> A_IWL<26632> A_IWL<26631> A_IWL<26630> A_IWL<26629> A_IWL<26628> A_IWL<26627> A_IWL<26626> A_IWL<26625> A_IWL<26624> A_IWL<27647> A_IWL<27646> A_IWL<27645> A_IWL<27644> A_IWL<27643> A_IWL<27642> A_IWL<27641> A_IWL<27640> A_IWL<27639> A_IWL<27638> A_IWL<27637> A_IWL<27636> A_IWL<27635> A_IWL<27634> A_IWL<27633> A_IWL<27632> A_IWL<27631> A_IWL<27630> A_IWL<27629> A_IWL<27628> A_IWL<27627> A_IWL<27626> A_IWL<27625> A_IWL<27624> A_IWL<27623> A_IWL<27622> A_IWL<27621> A_IWL<27620> A_IWL<27619> A_IWL<27618> A_IWL<27617> A_IWL<27616> A_IWL<27615> A_IWL<27614> A_IWL<27613> A_IWL<27612> A_IWL<27611> A_IWL<27610> A_IWL<27609> A_IWL<27608> A_IWL<27607> A_IWL<27606> A_IWL<27605> A_IWL<27604> A_IWL<27603> A_IWL<27602> A_IWL<27601> A_IWL<27600> A_IWL<27599> A_IWL<27598> A_IWL<27597> A_IWL<27596> A_IWL<27595> A_IWL<27594> A_IWL<27593> A_IWL<27592> A_IWL<27591> A_IWL<27590> A_IWL<27589> A_IWL<27588> A_IWL<27587> A_IWL<27586> A_IWL<27585> A_IWL<27584> A_IWL<27583> A_IWL<27582> A_IWL<27581> A_IWL<27580> A_IWL<27579> A_IWL<27578> A_IWL<27577> A_IWL<27576> A_IWL<27575> A_IWL<27574> A_IWL<27573> A_IWL<27572> A_IWL<27571> A_IWL<27570> A_IWL<27569> A_IWL<27568> A_IWL<27567> A_IWL<27566> A_IWL<27565> A_IWL<27564> A_IWL<27563> A_IWL<27562> A_IWL<27561> A_IWL<27560> A_IWL<27559> A_IWL<27558> A_IWL<27557> A_IWL<27556> A_IWL<27555> A_IWL<27554> A_IWL<27553> A_IWL<27552> A_IWL<27551> A_IWL<27550> A_IWL<27549> A_IWL<27548> A_IWL<27547> A_IWL<27546> A_IWL<27545> A_IWL<27544> A_IWL<27543> A_IWL<27542> A_IWL<27541> A_IWL<27540> A_IWL<27539> A_IWL<27538> A_IWL<27537> A_IWL<27536> A_IWL<27535> A_IWL<27534> A_IWL<27533> A_IWL<27532> A_IWL<27531> A_IWL<27530> A_IWL<27529> A_IWL<27528> A_IWL<27527> A_IWL<27526> A_IWL<27525> A_IWL<27524> A_IWL<27523> A_IWL<27522> A_IWL<27521> A_IWL<27520> A_IWL<27519> A_IWL<27518> A_IWL<27517> A_IWL<27516> A_IWL<27515> A_IWL<27514> A_IWL<27513> A_IWL<27512> A_IWL<27511> A_IWL<27510> A_IWL<27509> A_IWL<27508> A_IWL<27507> A_IWL<27506> A_IWL<27505> A_IWL<27504> A_IWL<27503> A_IWL<27502> A_IWL<27501> A_IWL<27500> A_IWL<27499> A_IWL<27498> A_IWL<27497> A_IWL<27496> A_IWL<27495> A_IWL<27494> A_IWL<27493> A_IWL<27492> A_IWL<27491> A_IWL<27490> A_IWL<27489> A_IWL<27488> A_IWL<27487> A_IWL<27486> A_IWL<27485> A_IWL<27484> A_IWL<27483> A_IWL<27482> A_IWL<27481> A_IWL<27480> A_IWL<27479> A_IWL<27478> A_IWL<27477> A_IWL<27476> A_IWL<27475> A_IWL<27474> A_IWL<27473> A_IWL<27472> A_IWL<27471> A_IWL<27470> A_IWL<27469> A_IWL<27468> A_IWL<27467> A_IWL<27466> A_IWL<27465> A_IWL<27464> A_IWL<27463> A_IWL<27462> A_IWL<27461> A_IWL<27460> A_IWL<27459> A_IWL<27458> A_IWL<27457> A_IWL<27456> A_IWL<27455> A_IWL<27454> A_IWL<27453> A_IWL<27452> A_IWL<27451> A_IWL<27450> A_IWL<27449> A_IWL<27448> A_IWL<27447> A_IWL<27446> A_IWL<27445> A_IWL<27444> A_IWL<27443> A_IWL<27442> A_IWL<27441> A_IWL<27440> A_IWL<27439> A_IWL<27438> A_IWL<27437> A_IWL<27436> A_IWL<27435> A_IWL<27434> A_IWL<27433> A_IWL<27432> A_IWL<27431> A_IWL<27430> A_IWL<27429> A_IWL<27428> A_IWL<27427> A_IWL<27426> A_IWL<27425> A_IWL<27424> A_IWL<27423> A_IWL<27422> A_IWL<27421> A_IWL<27420> A_IWL<27419> A_IWL<27418> A_IWL<27417> A_IWL<27416> A_IWL<27415> A_IWL<27414> A_IWL<27413> A_IWL<27412> A_IWL<27411> A_IWL<27410> A_IWL<27409> A_IWL<27408> A_IWL<27407> A_IWL<27406> A_IWL<27405> A_IWL<27404> A_IWL<27403> A_IWL<27402> A_IWL<27401> A_IWL<27400> A_IWL<27399> A_IWL<27398> A_IWL<27397> A_IWL<27396> A_IWL<27395> A_IWL<27394> A_IWL<27393> A_IWL<27392> A_IWL<27391> A_IWL<27390> A_IWL<27389> A_IWL<27388> A_IWL<27387> A_IWL<27386> A_IWL<27385> A_IWL<27384> A_IWL<27383> A_IWL<27382> A_IWL<27381> A_IWL<27380> A_IWL<27379> A_IWL<27378> A_IWL<27377> A_IWL<27376> A_IWL<27375> A_IWL<27374> A_IWL<27373> A_IWL<27372> A_IWL<27371> A_IWL<27370> A_IWL<27369> A_IWL<27368> A_IWL<27367> A_IWL<27366> A_IWL<27365> A_IWL<27364> A_IWL<27363> A_IWL<27362> A_IWL<27361> A_IWL<27360> A_IWL<27359> A_IWL<27358> A_IWL<27357> A_IWL<27356> A_IWL<27355> A_IWL<27354> A_IWL<27353> A_IWL<27352> A_IWL<27351> A_IWL<27350> A_IWL<27349> A_IWL<27348> A_IWL<27347> A_IWL<27346> A_IWL<27345> A_IWL<27344> A_IWL<27343> A_IWL<27342> A_IWL<27341> A_IWL<27340> A_IWL<27339> A_IWL<27338> A_IWL<27337> A_IWL<27336> A_IWL<27335> A_IWL<27334> A_IWL<27333> A_IWL<27332> A_IWL<27331> A_IWL<27330> A_IWL<27329> A_IWL<27328> A_IWL<27327> A_IWL<27326> A_IWL<27325> A_IWL<27324> A_IWL<27323> A_IWL<27322> A_IWL<27321> A_IWL<27320> A_IWL<27319> A_IWL<27318> A_IWL<27317> A_IWL<27316> A_IWL<27315> A_IWL<27314> A_IWL<27313> A_IWL<27312> A_IWL<27311> A_IWL<27310> A_IWL<27309> A_IWL<27308> A_IWL<27307> A_IWL<27306> A_IWL<27305> A_IWL<27304> A_IWL<27303> A_IWL<27302> A_IWL<27301> A_IWL<27300> A_IWL<27299> A_IWL<27298> A_IWL<27297> A_IWL<27296> A_IWL<27295> A_IWL<27294> A_IWL<27293> A_IWL<27292> A_IWL<27291> A_IWL<27290> A_IWL<27289> A_IWL<27288> A_IWL<27287> A_IWL<27286> A_IWL<27285> A_IWL<27284> A_IWL<27283> A_IWL<27282> A_IWL<27281> A_IWL<27280> A_IWL<27279> A_IWL<27278> A_IWL<27277> A_IWL<27276> A_IWL<27275> A_IWL<27274> A_IWL<27273> A_IWL<27272> A_IWL<27271> A_IWL<27270> A_IWL<27269> A_IWL<27268> A_IWL<27267> A_IWL<27266> A_IWL<27265> A_IWL<27264> A_IWL<27263> A_IWL<27262> A_IWL<27261> A_IWL<27260> A_IWL<27259> A_IWL<27258> A_IWL<27257> A_IWL<27256> A_IWL<27255> A_IWL<27254> A_IWL<27253> A_IWL<27252> A_IWL<27251> A_IWL<27250> A_IWL<27249> A_IWL<27248> A_IWL<27247> A_IWL<27246> A_IWL<27245> A_IWL<27244> A_IWL<27243> A_IWL<27242> A_IWL<27241> A_IWL<27240> A_IWL<27239> A_IWL<27238> A_IWL<27237> A_IWL<27236> A_IWL<27235> A_IWL<27234> A_IWL<27233> A_IWL<27232> A_IWL<27231> A_IWL<27230> A_IWL<27229> A_IWL<27228> A_IWL<27227> A_IWL<27226> A_IWL<27225> A_IWL<27224> A_IWL<27223> A_IWL<27222> A_IWL<27221> A_IWL<27220> A_IWL<27219> A_IWL<27218> A_IWL<27217> A_IWL<27216> A_IWL<27215> A_IWL<27214> A_IWL<27213> A_IWL<27212> A_IWL<27211> A_IWL<27210> A_IWL<27209> A_IWL<27208> A_IWL<27207> A_IWL<27206> A_IWL<27205> A_IWL<27204> A_IWL<27203> A_IWL<27202> A_IWL<27201> A_IWL<27200> A_IWL<27199> A_IWL<27198> A_IWL<27197> A_IWL<27196> A_IWL<27195> A_IWL<27194> A_IWL<27193> A_IWL<27192> A_IWL<27191> A_IWL<27190> A_IWL<27189> A_IWL<27188> A_IWL<27187> A_IWL<27186> A_IWL<27185> A_IWL<27184> A_IWL<27183> A_IWL<27182> A_IWL<27181> A_IWL<27180> A_IWL<27179> A_IWL<27178> A_IWL<27177> A_IWL<27176> A_IWL<27175> A_IWL<27174> A_IWL<27173> A_IWL<27172> A_IWL<27171> A_IWL<27170> A_IWL<27169> A_IWL<27168> A_IWL<27167> A_IWL<27166> A_IWL<27165> A_IWL<27164> A_IWL<27163> A_IWL<27162> A_IWL<27161> A_IWL<27160> A_IWL<27159> A_IWL<27158> A_IWL<27157> A_IWL<27156> A_IWL<27155> A_IWL<27154> A_IWL<27153> A_IWL<27152> A_IWL<27151> A_IWL<27150> A_IWL<27149> A_IWL<27148> A_IWL<27147> A_IWL<27146> A_IWL<27145> A_IWL<27144> A_IWL<27143> A_IWL<27142> A_IWL<27141> A_IWL<27140> A_IWL<27139> A_IWL<27138> A_IWL<27137> A_IWL<27136> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<52> A_BLC<105> A_BLC<104> A_BLC_TOP<105> A_BLC_TOP<104> A_BLT<105> A_BLT<104> A_BLT_TOP<105> A_BLT_TOP<104> A_IWL<26623> A_IWL<26622> A_IWL<26621> A_IWL<26620> A_IWL<26619> A_IWL<26618> A_IWL<26617> A_IWL<26616> A_IWL<26615> A_IWL<26614> A_IWL<26613> A_IWL<26612> A_IWL<26611> A_IWL<26610> A_IWL<26609> A_IWL<26608> A_IWL<26607> A_IWL<26606> A_IWL<26605> A_IWL<26604> A_IWL<26603> A_IWL<26602> A_IWL<26601> A_IWL<26600> A_IWL<26599> A_IWL<26598> A_IWL<26597> A_IWL<26596> A_IWL<26595> A_IWL<26594> A_IWL<26593> A_IWL<26592> A_IWL<26591> A_IWL<26590> A_IWL<26589> A_IWL<26588> A_IWL<26587> A_IWL<26586> A_IWL<26585> A_IWL<26584> A_IWL<26583> A_IWL<26582> A_IWL<26581> A_IWL<26580> A_IWL<26579> A_IWL<26578> A_IWL<26577> A_IWL<26576> A_IWL<26575> A_IWL<26574> A_IWL<26573> A_IWL<26572> A_IWL<26571> A_IWL<26570> A_IWL<26569> A_IWL<26568> A_IWL<26567> A_IWL<26566> A_IWL<26565> A_IWL<26564> A_IWL<26563> A_IWL<26562> A_IWL<26561> A_IWL<26560> A_IWL<26559> A_IWL<26558> A_IWL<26557> A_IWL<26556> A_IWL<26555> A_IWL<26554> A_IWL<26553> A_IWL<26552> A_IWL<26551> A_IWL<26550> A_IWL<26549> A_IWL<26548> A_IWL<26547> A_IWL<26546> A_IWL<26545> A_IWL<26544> A_IWL<26543> A_IWL<26542> A_IWL<26541> A_IWL<26540> A_IWL<26539> A_IWL<26538> A_IWL<26537> A_IWL<26536> A_IWL<26535> A_IWL<26534> A_IWL<26533> A_IWL<26532> A_IWL<26531> A_IWL<26530> A_IWL<26529> A_IWL<26528> A_IWL<26527> A_IWL<26526> A_IWL<26525> A_IWL<26524> A_IWL<26523> A_IWL<26522> A_IWL<26521> A_IWL<26520> A_IWL<26519> A_IWL<26518> A_IWL<26517> A_IWL<26516> A_IWL<26515> A_IWL<26514> A_IWL<26513> A_IWL<26512> A_IWL<26511> A_IWL<26510> A_IWL<26509> A_IWL<26508> A_IWL<26507> A_IWL<26506> A_IWL<26505> A_IWL<26504> A_IWL<26503> A_IWL<26502> A_IWL<26501> A_IWL<26500> A_IWL<26499> A_IWL<26498> A_IWL<26497> A_IWL<26496> A_IWL<26495> A_IWL<26494> A_IWL<26493> A_IWL<26492> A_IWL<26491> A_IWL<26490> A_IWL<26489> A_IWL<26488> A_IWL<26487> A_IWL<26486> A_IWL<26485> A_IWL<26484> A_IWL<26483> A_IWL<26482> A_IWL<26481> A_IWL<26480> A_IWL<26479> A_IWL<26478> A_IWL<26477> A_IWL<26476> A_IWL<26475> A_IWL<26474> A_IWL<26473> A_IWL<26472> A_IWL<26471> A_IWL<26470> A_IWL<26469> A_IWL<26468> A_IWL<26467> A_IWL<26466> A_IWL<26465> A_IWL<26464> A_IWL<26463> A_IWL<26462> A_IWL<26461> A_IWL<26460> A_IWL<26459> A_IWL<26458> A_IWL<26457> A_IWL<26456> A_IWL<26455> A_IWL<26454> A_IWL<26453> A_IWL<26452> A_IWL<26451> A_IWL<26450> A_IWL<26449> A_IWL<26448> A_IWL<26447> A_IWL<26446> A_IWL<26445> A_IWL<26444> A_IWL<26443> A_IWL<26442> A_IWL<26441> A_IWL<26440> A_IWL<26439> A_IWL<26438> A_IWL<26437> A_IWL<26436> A_IWL<26435> A_IWL<26434> A_IWL<26433> A_IWL<26432> A_IWL<26431> A_IWL<26430> A_IWL<26429> A_IWL<26428> A_IWL<26427> A_IWL<26426> A_IWL<26425> A_IWL<26424> A_IWL<26423> A_IWL<26422> A_IWL<26421> A_IWL<26420> A_IWL<26419> A_IWL<26418> A_IWL<26417> A_IWL<26416> A_IWL<26415> A_IWL<26414> A_IWL<26413> A_IWL<26412> A_IWL<26411> A_IWL<26410> A_IWL<26409> A_IWL<26408> A_IWL<26407> A_IWL<26406> A_IWL<26405> A_IWL<26404> A_IWL<26403> A_IWL<26402> A_IWL<26401> A_IWL<26400> A_IWL<26399> A_IWL<26398> A_IWL<26397> A_IWL<26396> A_IWL<26395> A_IWL<26394> A_IWL<26393> A_IWL<26392> A_IWL<26391> A_IWL<26390> A_IWL<26389> A_IWL<26388> A_IWL<26387> A_IWL<26386> A_IWL<26385> A_IWL<26384> A_IWL<26383> A_IWL<26382> A_IWL<26381> A_IWL<26380> A_IWL<26379> A_IWL<26378> A_IWL<26377> A_IWL<26376> A_IWL<26375> A_IWL<26374> A_IWL<26373> A_IWL<26372> A_IWL<26371> A_IWL<26370> A_IWL<26369> A_IWL<26368> A_IWL<26367> A_IWL<26366> A_IWL<26365> A_IWL<26364> A_IWL<26363> A_IWL<26362> A_IWL<26361> A_IWL<26360> A_IWL<26359> A_IWL<26358> A_IWL<26357> A_IWL<26356> A_IWL<26355> A_IWL<26354> A_IWL<26353> A_IWL<26352> A_IWL<26351> A_IWL<26350> A_IWL<26349> A_IWL<26348> A_IWL<26347> A_IWL<26346> A_IWL<26345> A_IWL<26344> A_IWL<26343> A_IWL<26342> A_IWL<26341> A_IWL<26340> A_IWL<26339> A_IWL<26338> A_IWL<26337> A_IWL<26336> A_IWL<26335> A_IWL<26334> A_IWL<26333> A_IWL<26332> A_IWL<26331> A_IWL<26330> A_IWL<26329> A_IWL<26328> A_IWL<26327> A_IWL<26326> A_IWL<26325> A_IWL<26324> A_IWL<26323> A_IWL<26322> A_IWL<26321> A_IWL<26320> A_IWL<26319> A_IWL<26318> A_IWL<26317> A_IWL<26316> A_IWL<26315> A_IWL<26314> A_IWL<26313> A_IWL<26312> A_IWL<26311> A_IWL<26310> A_IWL<26309> A_IWL<26308> A_IWL<26307> A_IWL<26306> A_IWL<26305> A_IWL<26304> A_IWL<26303> A_IWL<26302> A_IWL<26301> A_IWL<26300> A_IWL<26299> A_IWL<26298> A_IWL<26297> A_IWL<26296> A_IWL<26295> A_IWL<26294> A_IWL<26293> A_IWL<26292> A_IWL<26291> A_IWL<26290> A_IWL<26289> A_IWL<26288> A_IWL<26287> A_IWL<26286> A_IWL<26285> A_IWL<26284> A_IWL<26283> A_IWL<26282> A_IWL<26281> A_IWL<26280> A_IWL<26279> A_IWL<26278> A_IWL<26277> A_IWL<26276> A_IWL<26275> A_IWL<26274> A_IWL<26273> A_IWL<26272> A_IWL<26271> A_IWL<26270> A_IWL<26269> A_IWL<26268> A_IWL<26267> A_IWL<26266> A_IWL<26265> A_IWL<26264> A_IWL<26263> A_IWL<26262> A_IWL<26261> A_IWL<26260> A_IWL<26259> A_IWL<26258> A_IWL<26257> A_IWL<26256> A_IWL<26255> A_IWL<26254> A_IWL<26253> A_IWL<26252> A_IWL<26251> A_IWL<26250> A_IWL<26249> A_IWL<26248> A_IWL<26247> A_IWL<26246> A_IWL<26245> A_IWL<26244> A_IWL<26243> A_IWL<26242> A_IWL<26241> A_IWL<26240> A_IWL<26239> A_IWL<26238> A_IWL<26237> A_IWL<26236> A_IWL<26235> A_IWL<26234> A_IWL<26233> A_IWL<26232> A_IWL<26231> A_IWL<26230> A_IWL<26229> A_IWL<26228> A_IWL<26227> A_IWL<26226> A_IWL<26225> A_IWL<26224> A_IWL<26223> A_IWL<26222> A_IWL<26221> A_IWL<26220> A_IWL<26219> A_IWL<26218> A_IWL<26217> A_IWL<26216> A_IWL<26215> A_IWL<26214> A_IWL<26213> A_IWL<26212> A_IWL<26211> A_IWL<26210> A_IWL<26209> A_IWL<26208> A_IWL<26207> A_IWL<26206> A_IWL<26205> A_IWL<26204> A_IWL<26203> A_IWL<26202> A_IWL<26201> A_IWL<26200> A_IWL<26199> A_IWL<26198> A_IWL<26197> A_IWL<26196> A_IWL<26195> A_IWL<26194> A_IWL<26193> A_IWL<26192> A_IWL<26191> A_IWL<26190> A_IWL<26189> A_IWL<26188> A_IWL<26187> A_IWL<26186> A_IWL<26185> A_IWL<26184> A_IWL<26183> A_IWL<26182> A_IWL<26181> A_IWL<26180> A_IWL<26179> A_IWL<26178> A_IWL<26177> A_IWL<26176> A_IWL<26175> A_IWL<26174> A_IWL<26173> A_IWL<26172> A_IWL<26171> A_IWL<26170> A_IWL<26169> A_IWL<26168> A_IWL<26167> A_IWL<26166> A_IWL<26165> A_IWL<26164> A_IWL<26163> A_IWL<26162> A_IWL<26161> A_IWL<26160> A_IWL<26159> A_IWL<26158> A_IWL<26157> A_IWL<26156> A_IWL<26155> A_IWL<26154> A_IWL<26153> A_IWL<26152> A_IWL<26151> A_IWL<26150> A_IWL<26149> A_IWL<26148> A_IWL<26147> A_IWL<26146> A_IWL<26145> A_IWL<26144> A_IWL<26143> A_IWL<26142> A_IWL<26141> A_IWL<26140> A_IWL<26139> A_IWL<26138> A_IWL<26137> A_IWL<26136> A_IWL<26135> A_IWL<26134> A_IWL<26133> A_IWL<26132> A_IWL<26131> A_IWL<26130> A_IWL<26129> A_IWL<26128> A_IWL<26127> A_IWL<26126> A_IWL<26125> A_IWL<26124> A_IWL<26123> A_IWL<26122> A_IWL<26121> A_IWL<26120> A_IWL<26119> A_IWL<26118> A_IWL<26117> A_IWL<26116> A_IWL<26115> A_IWL<26114> A_IWL<26113> A_IWL<26112> A_IWL<27135> A_IWL<27134> A_IWL<27133> A_IWL<27132> A_IWL<27131> A_IWL<27130> A_IWL<27129> A_IWL<27128> A_IWL<27127> A_IWL<27126> A_IWL<27125> A_IWL<27124> A_IWL<27123> A_IWL<27122> A_IWL<27121> A_IWL<27120> A_IWL<27119> A_IWL<27118> A_IWL<27117> A_IWL<27116> A_IWL<27115> A_IWL<27114> A_IWL<27113> A_IWL<27112> A_IWL<27111> A_IWL<27110> A_IWL<27109> A_IWL<27108> A_IWL<27107> A_IWL<27106> A_IWL<27105> A_IWL<27104> A_IWL<27103> A_IWL<27102> A_IWL<27101> A_IWL<27100> A_IWL<27099> A_IWL<27098> A_IWL<27097> A_IWL<27096> A_IWL<27095> A_IWL<27094> A_IWL<27093> A_IWL<27092> A_IWL<27091> A_IWL<27090> A_IWL<27089> A_IWL<27088> A_IWL<27087> A_IWL<27086> A_IWL<27085> A_IWL<27084> A_IWL<27083> A_IWL<27082> A_IWL<27081> A_IWL<27080> A_IWL<27079> A_IWL<27078> A_IWL<27077> A_IWL<27076> A_IWL<27075> A_IWL<27074> A_IWL<27073> A_IWL<27072> A_IWL<27071> A_IWL<27070> A_IWL<27069> A_IWL<27068> A_IWL<27067> A_IWL<27066> A_IWL<27065> A_IWL<27064> A_IWL<27063> A_IWL<27062> A_IWL<27061> A_IWL<27060> A_IWL<27059> A_IWL<27058> A_IWL<27057> A_IWL<27056> A_IWL<27055> A_IWL<27054> A_IWL<27053> A_IWL<27052> A_IWL<27051> A_IWL<27050> A_IWL<27049> A_IWL<27048> A_IWL<27047> A_IWL<27046> A_IWL<27045> A_IWL<27044> A_IWL<27043> A_IWL<27042> A_IWL<27041> A_IWL<27040> A_IWL<27039> A_IWL<27038> A_IWL<27037> A_IWL<27036> A_IWL<27035> A_IWL<27034> A_IWL<27033> A_IWL<27032> A_IWL<27031> A_IWL<27030> A_IWL<27029> A_IWL<27028> A_IWL<27027> A_IWL<27026> A_IWL<27025> A_IWL<27024> A_IWL<27023> A_IWL<27022> A_IWL<27021> A_IWL<27020> A_IWL<27019> A_IWL<27018> A_IWL<27017> A_IWL<27016> A_IWL<27015> A_IWL<27014> A_IWL<27013> A_IWL<27012> A_IWL<27011> A_IWL<27010> A_IWL<27009> A_IWL<27008> A_IWL<27007> A_IWL<27006> A_IWL<27005> A_IWL<27004> A_IWL<27003> A_IWL<27002> A_IWL<27001> A_IWL<27000> A_IWL<26999> A_IWL<26998> A_IWL<26997> A_IWL<26996> A_IWL<26995> A_IWL<26994> A_IWL<26993> A_IWL<26992> A_IWL<26991> A_IWL<26990> A_IWL<26989> A_IWL<26988> A_IWL<26987> A_IWL<26986> A_IWL<26985> A_IWL<26984> A_IWL<26983> A_IWL<26982> A_IWL<26981> A_IWL<26980> A_IWL<26979> A_IWL<26978> A_IWL<26977> A_IWL<26976> A_IWL<26975> A_IWL<26974> A_IWL<26973> A_IWL<26972> A_IWL<26971> A_IWL<26970> A_IWL<26969> A_IWL<26968> A_IWL<26967> A_IWL<26966> A_IWL<26965> A_IWL<26964> A_IWL<26963> A_IWL<26962> A_IWL<26961> A_IWL<26960> A_IWL<26959> A_IWL<26958> A_IWL<26957> A_IWL<26956> A_IWL<26955> A_IWL<26954> A_IWL<26953> A_IWL<26952> A_IWL<26951> A_IWL<26950> A_IWL<26949> A_IWL<26948> A_IWL<26947> A_IWL<26946> A_IWL<26945> A_IWL<26944> A_IWL<26943> A_IWL<26942> A_IWL<26941> A_IWL<26940> A_IWL<26939> A_IWL<26938> A_IWL<26937> A_IWL<26936> A_IWL<26935> A_IWL<26934> A_IWL<26933> A_IWL<26932> A_IWL<26931> A_IWL<26930> A_IWL<26929> A_IWL<26928> A_IWL<26927> A_IWL<26926> A_IWL<26925> A_IWL<26924> A_IWL<26923> A_IWL<26922> A_IWL<26921> A_IWL<26920> A_IWL<26919> A_IWL<26918> A_IWL<26917> A_IWL<26916> A_IWL<26915> A_IWL<26914> A_IWL<26913> A_IWL<26912> A_IWL<26911> A_IWL<26910> A_IWL<26909> A_IWL<26908> A_IWL<26907> A_IWL<26906> A_IWL<26905> A_IWL<26904> A_IWL<26903> A_IWL<26902> A_IWL<26901> A_IWL<26900> A_IWL<26899> A_IWL<26898> A_IWL<26897> A_IWL<26896> A_IWL<26895> A_IWL<26894> A_IWL<26893> A_IWL<26892> A_IWL<26891> A_IWL<26890> A_IWL<26889> A_IWL<26888> A_IWL<26887> A_IWL<26886> A_IWL<26885> A_IWL<26884> A_IWL<26883> A_IWL<26882> A_IWL<26881> A_IWL<26880> A_IWL<26879> A_IWL<26878> A_IWL<26877> A_IWL<26876> A_IWL<26875> A_IWL<26874> A_IWL<26873> A_IWL<26872> A_IWL<26871> A_IWL<26870> A_IWL<26869> A_IWL<26868> A_IWL<26867> A_IWL<26866> A_IWL<26865> A_IWL<26864> A_IWL<26863> A_IWL<26862> A_IWL<26861> A_IWL<26860> A_IWL<26859> A_IWL<26858> A_IWL<26857> A_IWL<26856> A_IWL<26855> A_IWL<26854> A_IWL<26853> A_IWL<26852> A_IWL<26851> A_IWL<26850> A_IWL<26849> A_IWL<26848> A_IWL<26847> A_IWL<26846> A_IWL<26845> A_IWL<26844> A_IWL<26843> A_IWL<26842> A_IWL<26841> A_IWL<26840> A_IWL<26839> A_IWL<26838> A_IWL<26837> A_IWL<26836> A_IWL<26835> A_IWL<26834> A_IWL<26833> A_IWL<26832> A_IWL<26831> A_IWL<26830> A_IWL<26829> A_IWL<26828> A_IWL<26827> A_IWL<26826> A_IWL<26825> A_IWL<26824> A_IWL<26823> A_IWL<26822> A_IWL<26821> A_IWL<26820> A_IWL<26819> A_IWL<26818> A_IWL<26817> A_IWL<26816> A_IWL<26815> A_IWL<26814> A_IWL<26813> A_IWL<26812> A_IWL<26811> A_IWL<26810> A_IWL<26809> A_IWL<26808> A_IWL<26807> A_IWL<26806> A_IWL<26805> A_IWL<26804> A_IWL<26803> A_IWL<26802> A_IWL<26801> A_IWL<26800> A_IWL<26799> A_IWL<26798> A_IWL<26797> A_IWL<26796> A_IWL<26795> A_IWL<26794> A_IWL<26793> A_IWL<26792> A_IWL<26791> A_IWL<26790> A_IWL<26789> A_IWL<26788> A_IWL<26787> A_IWL<26786> A_IWL<26785> A_IWL<26784> A_IWL<26783> A_IWL<26782> A_IWL<26781> A_IWL<26780> A_IWL<26779> A_IWL<26778> A_IWL<26777> A_IWL<26776> A_IWL<26775> A_IWL<26774> A_IWL<26773> A_IWL<26772> A_IWL<26771> A_IWL<26770> A_IWL<26769> A_IWL<26768> A_IWL<26767> A_IWL<26766> A_IWL<26765> A_IWL<26764> A_IWL<26763> A_IWL<26762> A_IWL<26761> A_IWL<26760> A_IWL<26759> A_IWL<26758> A_IWL<26757> A_IWL<26756> A_IWL<26755> A_IWL<26754> A_IWL<26753> A_IWL<26752> A_IWL<26751> A_IWL<26750> A_IWL<26749> A_IWL<26748> A_IWL<26747> A_IWL<26746> A_IWL<26745> A_IWL<26744> A_IWL<26743> A_IWL<26742> A_IWL<26741> A_IWL<26740> A_IWL<26739> A_IWL<26738> A_IWL<26737> A_IWL<26736> A_IWL<26735> A_IWL<26734> A_IWL<26733> A_IWL<26732> A_IWL<26731> A_IWL<26730> A_IWL<26729> A_IWL<26728> A_IWL<26727> A_IWL<26726> A_IWL<26725> A_IWL<26724> A_IWL<26723> A_IWL<26722> A_IWL<26721> A_IWL<26720> A_IWL<26719> A_IWL<26718> A_IWL<26717> A_IWL<26716> A_IWL<26715> A_IWL<26714> A_IWL<26713> A_IWL<26712> A_IWL<26711> A_IWL<26710> A_IWL<26709> A_IWL<26708> A_IWL<26707> A_IWL<26706> A_IWL<26705> A_IWL<26704> A_IWL<26703> A_IWL<26702> A_IWL<26701> A_IWL<26700> A_IWL<26699> A_IWL<26698> A_IWL<26697> A_IWL<26696> A_IWL<26695> A_IWL<26694> A_IWL<26693> A_IWL<26692> A_IWL<26691> A_IWL<26690> A_IWL<26689> A_IWL<26688> A_IWL<26687> A_IWL<26686> A_IWL<26685> A_IWL<26684> A_IWL<26683> A_IWL<26682> A_IWL<26681> A_IWL<26680> A_IWL<26679> A_IWL<26678> A_IWL<26677> A_IWL<26676> A_IWL<26675> A_IWL<26674> A_IWL<26673> A_IWL<26672> A_IWL<26671> A_IWL<26670> A_IWL<26669> A_IWL<26668> A_IWL<26667> A_IWL<26666> A_IWL<26665> A_IWL<26664> A_IWL<26663> A_IWL<26662> A_IWL<26661> A_IWL<26660> A_IWL<26659> A_IWL<26658> A_IWL<26657> A_IWL<26656> A_IWL<26655> A_IWL<26654> A_IWL<26653> A_IWL<26652> A_IWL<26651> A_IWL<26650> A_IWL<26649> A_IWL<26648> A_IWL<26647> A_IWL<26646> A_IWL<26645> A_IWL<26644> A_IWL<26643> A_IWL<26642> A_IWL<26641> A_IWL<26640> A_IWL<26639> A_IWL<26638> A_IWL<26637> A_IWL<26636> A_IWL<26635> A_IWL<26634> A_IWL<26633> A_IWL<26632> A_IWL<26631> A_IWL<26630> A_IWL<26629> A_IWL<26628> A_IWL<26627> A_IWL<26626> A_IWL<26625> A_IWL<26624> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<51> A_BLC<103> A_BLC<102> A_BLC_TOP<103> A_BLC_TOP<102> A_BLT<103> A_BLT<102> A_BLT_TOP<103> A_BLT_TOP<102> A_IWL<26111> A_IWL<26110> A_IWL<26109> A_IWL<26108> A_IWL<26107> A_IWL<26106> A_IWL<26105> A_IWL<26104> A_IWL<26103> A_IWL<26102> A_IWL<26101> A_IWL<26100> A_IWL<26099> A_IWL<26098> A_IWL<26097> A_IWL<26096> A_IWL<26095> A_IWL<26094> A_IWL<26093> A_IWL<26092> A_IWL<26091> A_IWL<26090> A_IWL<26089> A_IWL<26088> A_IWL<26087> A_IWL<26086> A_IWL<26085> A_IWL<26084> A_IWL<26083> A_IWL<26082> A_IWL<26081> A_IWL<26080> A_IWL<26079> A_IWL<26078> A_IWL<26077> A_IWL<26076> A_IWL<26075> A_IWL<26074> A_IWL<26073> A_IWL<26072> A_IWL<26071> A_IWL<26070> A_IWL<26069> A_IWL<26068> A_IWL<26067> A_IWL<26066> A_IWL<26065> A_IWL<26064> A_IWL<26063> A_IWL<26062> A_IWL<26061> A_IWL<26060> A_IWL<26059> A_IWL<26058> A_IWL<26057> A_IWL<26056> A_IWL<26055> A_IWL<26054> A_IWL<26053> A_IWL<26052> A_IWL<26051> A_IWL<26050> A_IWL<26049> A_IWL<26048> A_IWL<26047> A_IWL<26046> A_IWL<26045> A_IWL<26044> A_IWL<26043> A_IWL<26042> A_IWL<26041> A_IWL<26040> A_IWL<26039> A_IWL<26038> A_IWL<26037> A_IWL<26036> A_IWL<26035> A_IWL<26034> A_IWL<26033> A_IWL<26032> A_IWL<26031> A_IWL<26030> A_IWL<26029> A_IWL<26028> A_IWL<26027> A_IWL<26026> A_IWL<26025> A_IWL<26024> A_IWL<26023> A_IWL<26022> A_IWL<26021> A_IWL<26020> A_IWL<26019> A_IWL<26018> A_IWL<26017> A_IWL<26016> A_IWL<26015> A_IWL<26014> A_IWL<26013> A_IWL<26012> A_IWL<26011> A_IWL<26010> A_IWL<26009> A_IWL<26008> A_IWL<26007> A_IWL<26006> A_IWL<26005> A_IWL<26004> A_IWL<26003> A_IWL<26002> A_IWL<26001> A_IWL<26000> A_IWL<25999> A_IWL<25998> A_IWL<25997> A_IWL<25996> A_IWL<25995> A_IWL<25994> A_IWL<25993> A_IWL<25992> A_IWL<25991> A_IWL<25990> A_IWL<25989> A_IWL<25988> A_IWL<25987> A_IWL<25986> A_IWL<25985> A_IWL<25984> A_IWL<25983> A_IWL<25982> A_IWL<25981> A_IWL<25980> A_IWL<25979> A_IWL<25978> A_IWL<25977> A_IWL<25976> A_IWL<25975> A_IWL<25974> A_IWL<25973> A_IWL<25972> A_IWL<25971> A_IWL<25970> A_IWL<25969> A_IWL<25968> A_IWL<25967> A_IWL<25966> A_IWL<25965> A_IWL<25964> A_IWL<25963> A_IWL<25962> A_IWL<25961> A_IWL<25960> A_IWL<25959> A_IWL<25958> A_IWL<25957> A_IWL<25956> A_IWL<25955> A_IWL<25954> A_IWL<25953> A_IWL<25952> A_IWL<25951> A_IWL<25950> A_IWL<25949> A_IWL<25948> A_IWL<25947> A_IWL<25946> A_IWL<25945> A_IWL<25944> A_IWL<25943> A_IWL<25942> A_IWL<25941> A_IWL<25940> A_IWL<25939> A_IWL<25938> A_IWL<25937> A_IWL<25936> A_IWL<25935> A_IWL<25934> A_IWL<25933> A_IWL<25932> A_IWL<25931> A_IWL<25930> A_IWL<25929> A_IWL<25928> A_IWL<25927> A_IWL<25926> A_IWL<25925> A_IWL<25924> A_IWL<25923> A_IWL<25922> A_IWL<25921> A_IWL<25920> A_IWL<25919> A_IWL<25918> A_IWL<25917> A_IWL<25916> A_IWL<25915> A_IWL<25914> A_IWL<25913> A_IWL<25912> A_IWL<25911> A_IWL<25910> A_IWL<25909> A_IWL<25908> A_IWL<25907> A_IWL<25906> A_IWL<25905> A_IWL<25904> A_IWL<25903> A_IWL<25902> A_IWL<25901> A_IWL<25900> A_IWL<25899> A_IWL<25898> A_IWL<25897> A_IWL<25896> A_IWL<25895> A_IWL<25894> A_IWL<25893> A_IWL<25892> A_IWL<25891> A_IWL<25890> A_IWL<25889> A_IWL<25888> A_IWL<25887> A_IWL<25886> A_IWL<25885> A_IWL<25884> A_IWL<25883> A_IWL<25882> A_IWL<25881> A_IWL<25880> A_IWL<25879> A_IWL<25878> A_IWL<25877> A_IWL<25876> A_IWL<25875> A_IWL<25874> A_IWL<25873> A_IWL<25872> A_IWL<25871> A_IWL<25870> A_IWL<25869> A_IWL<25868> A_IWL<25867> A_IWL<25866> A_IWL<25865> A_IWL<25864> A_IWL<25863> A_IWL<25862> A_IWL<25861> A_IWL<25860> A_IWL<25859> A_IWL<25858> A_IWL<25857> A_IWL<25856> A_IWL<25855> A_IWL<25854> A_IWL<25853> A_IWL<25852> A_IWL<25851> A_IWL<25850> A_IWL<25849> A_IWL<25848> A_IWL<25847> A_IWL<25846> A_IWL<25845> A_IWL<25844> A_IWL<25843> A_IWL<25842> A_IWL<25841> A_IWL<25840> A_IWL<25839> A_IWL<25838> A_IWL<25837> A_IWL<25836> A_IWL<25835> A_IWL<25834> A_IWL<25833> A_IWL<25832> A_IWL<25831> A_IWL<25830> A_IWL<25829> A_IWL<25828> A_IWL<25827> A_IWL<25826> A_IWL<25825> A_IWL<25824> A_IWL<25823> A_IWL<25822> A_IWL<25821> A_IWL<25820> A_IWL<25819> A_IWL<25818> A_IWL<25817> A_IWL<25816> A_IWL<25815> A_IWL<25814> A_IWL<25813> A_IWL<25812> A_IWL<25811> A_IWL<25810> A_IWL<25809> A_IWL<25808> A_IWL<25807> A_IWL<25806> A_IWL<25805> A_IWL<25804> A_IWL<25803> A_IWL<25802> A_IWL<25801> A_IWL<25800> A_IWL<25799> A_IWL<25798> A_IWL<25797> A_IWL<25796> A_IWL<25795> A_IWL<25794> A_IWL<25793> A_IWL<25792> A_IWL<25791> A_IWL<25790> A_IWL<25789> A_IWL<25788> A_IWL<25787> A_IWL<25786> A_IWL<25785> A_IWL<25784> A_IWL<25783> A_IWL<25782> A_IWL<25781> A_IWL<25780> A_IWL<25779> A_IWL<25778> A_IWL<25777> A_IWL<25776> A_IWL<25775> A_IWL<25774> A_IWL<25773> A_IWL<25772> A_IWL<25771> A_IWL<25770> A_IWL<25769> A_IWL<25768> A_IWL<25767> A_IWL<25766> A_IWL<25765> A_IWL<25764> A_IWL<25763> A_IWL<25762> A_IWL<25761> A_IWL<25760> A_IWL<25759> A_IWL<25758> A_IWL<25757> A_IWL<25756> A_IWL<25755> A_IWL<25754> A_IWL<25753> A_IWL<25752> A_IWL<25751> A_IWL<25750> A_IWL<25749> A_IWL<25748> A_IWL<25747> A_IWL<25746> A_IWL<25745> A_IWL<25744> A_IWL<25743> A_IWL<25742> A_IWL<25741> A_IWL<25740> A_IWL<25739> A_IWL<25738> A_IWL<25737> A_IWL<25736> A_IWL<25735> A_IWL<25734> A_IWL<25733> A_IWL<25732> A_IWL<25731> A_IWL<25730> A_IWL<25729> A_IWL<25728> A_IWL<25727> A_IWL<25726> A_IWL<25725> A_IWL<25724> A_IWL<25723> A_IWL<25722> A_IWL<25721> A_IWL<25720> A_IWL<25719> A_IWL<25718> A_IWL<25717> A_IWL<25716> A_IWL<25715> A_IWL<25714> A_IWL<25713> A_IWL<25712> A_IWL<25711> A_IWL<25710> A_IWL<25709> A_IWL<25708> A_IWL<25707> A_IWL<25706> A_IWL<25705> A_IWL<25704> A_IWL<25703> A_IWL<25702> A_IWL<25701> A_IWL<25700> A_IWL<25699> A_IWL<25698> A_IWL<25697> A_IWL<25696> A_IWL<25695> A_IWL<25694> A_IWL<25693> A_IWL<25692> A_IWL<25691> A_IWL<25690> A_IWL<25689> A_IWL<25688> A_IWL<25687> A_IWL<25686> A_IWL<25685> A_IWL<25684> A_IWL<25683> A_IWL<25682> A_IWL<25681> A_IWL<25680> A_IWL<25679> A_IWL<25678> A_IWL<25677> A_IWL<25676> A_IWL<25675> A_IWL<25674> A_IWL<25673> A_IWL<25672> A_IWL<25671> A_IWL<25670> A_IWL<25669> A_IWL<25668> A_IWL<25667> A_IWL<25666> A_IWL<25665> A_IWL<25664> A_IWL<25663> A_IWL<25662> A_IWL<25661> A_IWL<25660> A_IWL<25659> A_IWL<25658> A_IWL<25657> A_IWL<25656> A_IWL<25655> A_IWL<25654> A_IWL<25653> A_IWL<25652> A_IWL<25651> A_IWL<25650> A_IWL<25649> A_IWL<25648> A_IWL<25647> A_IWL<25646> A_IWL<25645> A_IWL<25644> A_IWL<25643> A_IWL<25642> A_IWL<25641> A_IWL<25640> A_IWL<25639> A_IWL<25638> A_IWL<25637> A_IWL<25636> A_IWL<25635> A_IWL<25634> A_IWL<25633> A_IWL<25632> A_IWL<25631> A_IWL<25630> A_IWL<25629> A_IWL<25628> A_IWL<25627> A_IWL<25626> A_IWL<25625> A_IWL<25624> A_IWL<25623> A_IWL<25622> A_IWL<25621> A_IWL<25620> A_IWL<25619> A_IWL<25618> A_IWL<25617> A_IWL<25616> A_IWL<25615> A_IWL<25614> A_IWL<25613> A_IWL<25612> A_IWL<25611> A_IWL<25610> A_IWL<25609> A_IWL<25608> A_IWL<25607> A_IWL<25606> A_IWL<25605> A_IWL<25604> A_IWL<25603> A_IWL<25602> A_IWL<25601> A_IWL<25600> A_IWL<26623> A_IWL<26622> A_IWL<26621> A_IWL<26620> A_IWL<26619> A_IWL<26618> A_IWL<26617> A_IWL<26616> A_IWL<26615> A_IWL<26614> A_IWL<26613> A_IWL<26612> A_IWL<26611> A_IWL<26610> A_IWL<26609> A_IWL<26608> A_IWL<26607> A_IWL<26606> A_IWL<26605> A_IWL<26604> A_IWL<26603> A_IWL<26602> A_IWL<26601> A_IWL<26600> A_IWL<26599> A_IWL<26598> A_IWL<26597> A_IWL<26596> A_IWL<26595> A_IWL<26594> A_IWL<26593> A_IWL<26592> A_IWL<26591> A_IWL<26590> A_IWL<26589> A_IWL<26588> A_IWL<26587> A_IWL<26586> A_IWL<26585> A_IWL<26584> A_IWL<26583> A_IWL<26582> A_IWL<26581> A_IWL<26580> A_IWL<26579> A_IWL<26578> A_IWL<26577> A_IWL<26576> A_IWL<26575> A_IWL<26574> A_IWL<26573> A_IWL<26572> A_IWL<26571> A_IWL<26570> A_IWL<26569> A_IWL<26568> A_IWL<26567> A_IWL<26566> A_IWL<26565> A_IWL<26564> A_IWL<26563> A_IWL<26562> A_IWL<26561> A_IWL<26560> A_IWL<26559> A_IWL<26558> A_IWL<26557> A_IWL<26556> A_IWL<26555> A_IWL<26554> A_IWL<26553> A_IWL<26552> A_IWL<26551> A_IWL<26550> A_IWL<26549> A_IWL<26548> A_IWL<26547> A_IWL<26546> A_IWL<26545> A_IWL<26544> A_IWL<26543> A_IWL<26542> A_IWL<26541> A_IWL<26540> A_IWL<26539> A_IWL<26538> A_IWL<26537> A_IWL<26536> A_IWL<26535> A_IWL<26534> A_IWL<26533> A_IWL<26532> A_IWL<26531> A_IWL<26530> A_IWL<26529> A_IWL<26528> A_IWL<26527> A_IWL<26526> A_IWL<26525> A_IWL<26524> A_IWL<26523> A_IWL<26522> A_IWL<26521> A_IWL<26520> A_IWL<26519> A_IWL<26518> A_IWL<26517> A_IWL<26516> A_IWL<26515> A_IWL<26514> A_IWL<26513> A_IWL<26512> A_IWL<26511> A_IWL<26510> A_IWL<26509> A_IWL<26508> A_IWL<26507> A_IWL<26506> A_IWL<26505> A_IWL<26504> A_IWL<26503> A_IWL<26502> A_IWL<26501> A_IWL<26500> A_IWL<26499> A_IWL<26498> A_IWL<26497> A_IWL<26496> A_IWL<26495> A_IWL<26494> A_IWL<26493> A_IWL<26492> A_IWL<26491> A_IWL<26490> A_IWL<26489> A_IWL<26488> A_IWL<26487> A_IWL<26486> A_IWL<26485> A_IWL<26484> A_IWL<26483> A_IWL<26482> A_IWL<26481> A_IWL<26480> A_IWL<26479> A_IWL<26478> A_IWL<26477> A_IWL<26476> A_IWL<26475> A_IWL<26474> A_IWL<26473> A_IWL<26472> A_IWL<26471> A_IWL<26470> A_IWL<26469> A_IWL<26468> A_IWL<26467> A_IWL<26466> A_IWL<26465> A_IWL<26464> A_IWL<26463> A_IWL<26462> A_IWL<26461> A_IWL<26460> A_IWL<26459> A_IWL<26458> A_IWL<26457> A_IWL<26456> A_IWL<26455> A_IWL<26454> A_IWL<26453> A_IWL<26452> A_IWL<26451> A_IWL<26450> A_IWL<26449> A_IWL<26448> A_IWL<26447> A_IWL<26446> A_IWL<26445> A_IWL<26444> A_IWL<26443> A_IWL<26442> A_IWL<26441> A_IWL<26440> A_IWL<26439> A_IWL<26438> A_IWL<26437> A_IWL<26436> A_IWL<26435> A_IWL<26434> A_IWL<26433> A_IWL<26432> A_IWL<26431> A_IWL<26430> A_IWL<26429> A_IWL<26428> A_IWL<26427> A_IWL<26426> A_IWL<26425> A_IWL<26424> A_IWL<26423> A_IWL<26422> A_IWL<26421> A_IWL<26420> A_IWL<26419> A_IWL<26418> A_IWL<26417> A_IWL<26416> A_IWL<26415> A_IWL<26414> A_IWL<26413> A_IWL<26412> A_IWL<26411> A_IWL<26410> A_IWL<26409> A_IWL<26408> A_IWL<26407> A_IWL<26406> A_IWL<26405> A_IWL<26404> A_IWL<26403> A_IWL<26402> A_IWL<26401> A_IWL<26400> A_IWL<26399> A_IWL<26398> A_IWL<26397> A_IWL<26396> A_IWL<26395> A_IWL<26394> A_IWL<26393> A_IWL<26392> A_IWL<26391> A_IWL<26390> A_IWL<26389> A_IWL<26388> A_IWL<26387> A_IWL<26386> A_IWL<26385> A_IWL<26384> A_IWL<26383> A_IWL<26382> A_IWL<26381> A_IWL<26380> A_IWL<26379> A_IWL<26378> A_IWL<26377> A_IWL<26376> A_IWL<26375> A_IWL<26374> A_IWL<26373> A_IWL<26372> A_IWL<26371> A_IWL<26370> A_IWL<26369> A_IWL<26368> A_IWL<26367> A_IWL<26366> A_IWL<26365> A_IWL<26364> A_IWL<26363> A_IWL<26362> A_IWL<26361> A_IWL<26360> A_IWL<26359> A_IWL<26358> A_IWL<26357> A_IWL<26356> A_IWL<26355> A_IWL<26354> A_IWL<26353> A_IWL<26352> A_IWL<26351> A_IWL<26350> A_IWL<26349> A_IWL<26348> A_IWL<26347> A_IWL<26346> A_IWL<26345> A_IWL<26344> A_IWL<26343> A_IWL<26342> A_IWL<26341> A_IWL<26340> A_IWL<26339> A_IWL<26338> A_IWL<26337> A_IWL<26336> A_IWL<26335> A_IWL<26334> A_IWL<26333> A_IWL<26332> A_IWL<26331> A_IWL<26330> A_IWL<26329> A_IWL<26328> A_IWL<26327> A_IWL<26326> A_IWL<26325> A_IWL<26324> A_IWL<26323> A_IWL<26322> A_IWL<26321> A_IWL<26320> A_IWL<26319> A_IWL<26318> A_IWL<26317> A_IWL<26316> A_IWL<26315> A_IWL<26314> A_IWL<26313> A_IWL<26312> A_IWL<26311> A_IWL<26310> A_IWL<26309> A_IWL<26308> A_IWL<26307> A_IWL<26306> A_IWL<26305> A_IWL<26304> A_IWL<26303> A_IWL<26302> A_IWL<26301> A_IWL<26300> A_IWL<26299> A_IWL<26298> A_IWL<26297> A_IWL<26296> A_IWL<26295> A_IWL<26294> A_IWL<26293> A_IWL<26292> A_IWL<26291> A_IWL<26290> A_IWL<26289> A_IWL<26288> A_IWL<26287> A_IWL<26286> A_IWL<26285> A_IWL<26284> A_IWL<26283> A_IWL<26282> A_IWL<26281> A_IWL<26280> A_IWL<26279> A_IWL<26278> A_IWL<26277> A_IWL<26276> A_IWL<26275> A_IWL<26274> A_IWL<26273> A_IWL<26272> A_IWL<26271> A_IWL<26270> A_IWL<26269> A_IWL<26268> A_IWL<26267> A_IWL<26266> A_IWL<26265> A_IWL<26264> A_IWL<26263> A_IWL<26262> A_IWL<26261> A_IWL<26260> A_IWL<26259> A_IWL<26258> A_IWL<26257> A_IWL<26256> A_IWL<26255> A_IWL<26254> A_IWL<26253> A_IWL<26252> A_IWL<26251> A_IWL<26250> A_IWL<26249> A_IWL<26248> A_IWL<26247> A_IWL<26246> A_IWL<26245> A_IWL<26244> A_IWL<26243> A_IWL<26242> A_IWL<26241> A_IWL<26240> A_IWL<26239> A_IWL<26238> A_IWL<26237> A_IWL<26236> A_IWL<26235> A_IWL<26234> A_IWL<26233> A_IWL<26232> A_IWL<26231> A_IWL<26230> A_IWL<26229> A_IWL<26228> A_IWL<26227> A_IWL<26226> A_IWL<26225> A_IWL<26224> A_IWL<26223> A_IWL<26222> A_IWL<26221> A_IWL<26220> A_IWL<26219> A_IWL<26218> A_IWL<26217> A_IWL<26216> A_IWL<26215> A_IWL<26214> A_IWL<26213> A_IWL<26212> A_IWL<26211> A_IWL<26210> A_IWL<26209> A_IWL<26208> A_IWL<26207> A_IWL<26206> A_IWL<26205> A_IWL<26204> A_IWL<26203> A_IWL<26202> A_IWL<26201> A_IWL<26200> A_IWL<26199> A_IWL<26198> A_IWL<26197> A_IWL<26196> A_IWL<26195> A_IWL<26194> A_IWL<26193> A_IWL<26192> A_IWL<26191> A_IWL<26190> A_IWL<26189> A_IWL<26188> A_IWL<26187> A_IWL<26186> A_IWL<26185> A_IWL<26184> A_IWL<26183> A_IWL<26182> A_IWL<26181> A_IWL<26180> A_IWL<26179> A_IWL<26178> A_IWL<26177> A_IWL<26176> A_IWL<26175> A_IWL<26174> A_IWL<26173> A_IWL<26172> A_IWL<26171> A_IWL<26170> A_IWL<26169> A_IWL<26168> A_IWL<26167> A_IWL<26166> A_IWL<26165> A_IWL<26164> A_IWL<26163> A_IWL<26162> A_IWL<26161> A_IWL<26160> A_IWL<26159> A_IWL<26158> A_IWL<26157> A_IWL<26156> A_IWL<26155> A_IWL<26154> A_IWL<26153> A_IWL<26152> A_IWL<26151> A_IWL<26150> A_IWL<26149> A_IWL<26148> A_IWL<26147> A_IWL<26146> A_IWL<26145> A_IWL<26144> A_IWL<26143> A_IWL<26142> A_IWL<26141> A_IWL<26140> A_IWL<26139> A_IWL<26138> A_IWL<26137> A_IWL<26136> A_IWL<26135> A_IWL<26134> A_IWL<26133> A_IWL<26132> A_IWL<26131> A_IWL<26130> A_IWL<26129> A_IWL<26128> A_IWL<26127> A_IWL<26126> A_IWL<26125> A_IWL<26124> A_IWL<26123> A_IWL<26122> A_IWL<26121> A_IWL<26120> A_IWL<26119> A_IWL<26118> A_IWL<26117> A_IWL<26116> A_IWL<26115> A_IWL<26114> A_IWL<26113> A_IWL<26112> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<50> A_BLC<101> A_BLC<100> A_BLC_TOP<101> A_BLC_TOP<100> A_BLT<101> A_BLT<100> A_BLT_TOP<101> A_BLT_TOP<100> A_IWL<25599> A_IWL<25598> A_IWL<25597> A_IWL<25596> A_IWL<25595> A_IWL<25594> A_IWL<25593> A_IWL<25592> A_IWL<25591> A_IWL<25590> A_IWL<25589> A_IWL<25588> A_IWL<25587> A_IWL<25586> A_IWL<25585> A_IWL<25584> A_IWL<25583> A_IWL<25582> A_IWL<25581> A_IWL<25580> A_IWL<25579> A_IWL<25578> A_IWL<25577> A_IWL<25576> A_IWL<25575> A_IWL<25574> A_IWL<25573> A_IWL<25572> A_IWL<25571> A_IWL<25570> A_IWL<25569> A_IWL<25568> A_IWL<25567> A_IWL<25566> A_IWL<25565> A_IWL<25564> A_IWL<25563> A_IWL<25562> A_IWL<25561> A_IWL<25560> A_IWL<25559> A_IWL<25558> A_IWL<25557> A_IWL<25556> A_IWL<25555> A_IWL<25554> A_IWL<25553> A_IWL<25552> A_IWL<25551> A_IWL<25550> A_IWL<25549> A_IWL<25548> A_IWL<25547> A_IWL<25546> A_IWL<25545> A_IWL<25544> A_IWL<25543> A_IWL<25542> A_IWL<25541> A_IWL<25540> A_IWL<25539> A_IWL<25538> A_IWL<25537> A_IWL<25536> A_IWL<25535> A_IWL<25534> A_IWL<25533> A_IWL<25532> A_IWL<25531> A_IWL<25530> A_IWL<25529> A_IWL<25528> A_IWL<25527> A_IWL<25526> A_IWL<25525> A_IWL<25524> A_IWL<25523> A_IWL<25522> A_IWL<25521> A_IWL<25520> A_IWL<25519> A_IWL<25518> A_IWL<25517> A_IWL<25516> A_IWL<25515> A_IWL<25514> A_IWL<25513> A_IWL<25512> A_IWL<25511> A_IWL<25510> A_IWL<25509> A_IWL<25508> A_IWL<25507> A_IWL<25506> A_IWL<25505> A_IWL<25504> A_IWL<25503> A_IWL<25502> A_IWL<25501> A_IWL<25500> A_IWL<25499> A_IWL<25498> A_IWL<25497> A_IWL<25496> A_IWL<25495> A_IWL<25494> A_IWL<25493> A_IWL<25492> A_IWL<25491> A_IWL<25490> A_IWL<25489> A_IWL<25488> A_IWL<25487> A_IWL<25486> A_IWL<25485> A_IWL<25484> A_IWL<25483> A_IWL<25482> A_IWL<25481> A_IWL<25480> A_IWL<25479> A_IWL<25478> A_IWL<25477> A_IWL<25476> A_IWL<25475> A_IWL<25474> A_IWL<25473> A_IWL<25472> A_IWL<25471> A_IWL<25470> A_IWL<25469> A_IWL<25468> A_IWL<25467> A_IWL<25466> A_IWL<25465> A_IWL<25464> A_IWL<25463> A_IWL<25462> A_IWL<25461> A_IWL<25460> A_IWL<25459> A_IWL<25458> A_IWL<25457> A_IWL<25456> A_IWL<25455> A_IWL<25454> A_IWL<25453> A_IWL<25452> A_IWL<25451> A_IWL<25450> A_IWL<25449> A_IWL<25448> A_IWL<25447> A_IWL<25446> A_IWL<25445> A_IWL<25444> A_IWL<25443> A_IWL<25442> A_IWL<25441> A_IWL<25440> A_IWL<25439> A_IWL<25438> A_IWL<25437> A_IWL<25436> A_IWL<25435> A_IWL<25434> A_IWL<25433> A_IWL<25432> A_IWL<25431> A_IWL<25430> A_IWL<25429> A_IWL<25428> A_IWL<25427> A_IWL<25426> A_IWL<25425> A_IWL<25424> A_IWL<25423> A_IWL<25422> A_IWL<25421> A_IWL<25420> A_IWL<25419> A_IWL<25418> A_IWL<25417> A_IWL<25416> A_IWL<25415> A_IWL<25414> A_IWL<25413> A_IWL<25412> A_IWL<25411> A_IWL<25410> A_IWL<25409> A_IWL<25408> A_IWL<25407> A_IWL<25406> A_IWL<25405> A_IWL<25404> A_IWL<25403> A_IWL<25402> A_IWL<25401> A_IWL<25400> A_IWL<25399> A_IWL<25398> A_IWL<25397> A_IWL<25396> A_IWL<25395> A_IWL<25394> A_IWL<25393> A_IWL<25392> A_IWL<25391> A_IWL<25390> A_IWL<25389> A_IWL<25388> A_IWL<25387> A_IWL<25386> A_IWL<25385> A_IWL<25384> A_IWL<25383> A_IWL<25382> A_IWL<25381> A_IWL<25380> A_IWL<25379> A_IWL<25378> A_IWL<25377> A_IWL<25376> A_IWL<25375> A_IWL<25374> A_IWL<25373> A_IWL<25372> A_IWL<25371> A_IWL<25370> A_IWL<25369> A_IWL<25368> A_IWL<25367> A_IWL<25366> A_IWL<25365> A_IWL<25364> A_IWL<25363> A_IWL<25362> A_IWL<25361> A_IWL<25360> A_IWL<25359> A_IWL<25358> A_IWL<25357> A_IWL<25356> A_IWL<25355> A_IWL<25354> A_IWL<25353> A_IWL<25352> A_IWL<25351> A_IWL<25350> A_IWL<25349> A_IWL<25348> A_IWL<25347> A_IWL<25346> A_IWL<25345> A_IWL<25344> A_IWL<25343> A_IWL<25342> A_IWL<25341> A_IWL<25340> A_IWL<25339> A_IWL<25338> A_IWL<25337> A_IWL<25336> A_IWL<25335> A_IWL<25334> A_IWL<25333> A_IWL<25332> A_IWL<25331> A_IWL<25330> A_IWL<25329> A_IWL<25328> A_IWL<25327> A_IWL<25326> A_IWL<25325> A_IWL<25324> A_IWL<25323> A_IWL<25322> A_IWL<25321> A_IWL<25320> A_IWL<25319> A_IWL<25318> A_IWL<25317> A_IWL<25316> A_IWL<25315> A_IWL<25314> A_IWL<25313> A_IWL<25312> A_IWL<25311> A_IWL<25310> A_IWL<25309> A_IWL<25308> A_IWL<25307> A_IWL<25306> A_IWL<25305> A_IWL<25304> A_IWL<25303> A_IWL<25302> A_IWL<25301> A_IWL<25300> A_IWL<25299> A_IWL<25298> A_IWL<25297> A_IWL<25296> A_IWL<25295> A_IWL<25294> A_IWL<25293> A_IWL<25292> A_IWL<25291> A_IWL<25290> A_IWL<25289> A_IWL<25288> A_IWL<25287> A_IWL<25286> A_IWL<25285> A_IWL<25284> A_IWL<25283> A_IWL<25282> A_IWL<25281> A_IWL<25280> A_IWL<25279> A_IWL<25278> A_IWL<25277> A_IWL<25276> A_IWL<25275> A_IWL<25274> A_IWL<25273> A_IWL<25272> A_IWL<25271> A_IWL<25270> A_IWL<25269> A_IWL<25268> A_IWL<25267> A_IWL<25266> A_IWL<25265> A_IWL<25264> A_IWL<25263> A_IWL<25262> A_IWL<25261> A_IWL<25260> A_IWL<25259> A_IWL<25258> A_IWL<25257> A_IWL<25256> A_IWL<25255> A_IWL<25254> A_IWL<25253> A_IWL<25252> A_IWL<25251> A_IWL<25250> A_IWL<25249> A_IWL<25248> A_IWL<25247> A_IWL<25246> A_IWL<25245> A_IWL<25244> A_IWL<25243> A_IWL<25242> A_IWL<25241> A_IWL<25240> A_IWL<25239> A_IWL<25238> A_IWL<25237> A_IWL<25236> A_IWL<25235> A_IWL<25234> A_IWL<25233> A_IWL<25232> A_IWL<25231> A_IWL<25230> A_IWL<25229> A_IWL<25228> A_IWL<25227> A_IWL<25226> A_IWL<25225> A_IWL<25224> A_IWL<25223> A_IWL<25222> A_IWL<25221> A_IWL<25220> A_IWL<25219> A_IWL<25218> A_IWL<25217> A_IWL<25216> A_IWL<25215> A_IWL<25214> A_IWL<25213> A_IWL<25212> A_IWL<25211> A_IWL<25210> A_IWL<25209> A_IWL<25208> A_IWL<25207> A_IWL<25206> A_IWL<25205> A_IWL<25204> A_IWL<25203> A_IWL<25202> A_IWL<25201> A_IWL<25200> A_IWL<25199> A_IWL<25198> A_IWL<25197> A_IWL<25196> A_IWL<25195> A_IWL<25194> A_IWL<25193> A_IWL<25192> A_IWL<25191> A_IWL<25190> A_IWL<25189> A_IWL<25188> A_IWL<25187> A_IWL<25186> A_IWL<25185> A_IWL<25184> A_IWL<25183> A_IWL<25182> A_IWL<25181> A_IWL<25180> A_IWL<25179> A_IWL<25178> A_IWL<25177> A_IWL<25176> A_IWL<25175> A_IWL<25174> A_IWL<25173> A_IWL<25172> A_IWL<25171> A_IWL<25170> A_IWL<25169> A_IWL<25168> A_IWL<25167> A_IWL<25166> A_IWL<25165> A_IWL<25164> A_IWL<25163> A_IWL<25162> A_IWL<25161> A_IWL<25160> A_IWL<25159> A_IWL<25158> A_IWL<25157> A_IWL<25156> A_IWL<25155> A_IWL<25154> A_IWL<25153> A_IWL<25152> A_IWL<25151> A_IWL<25150> A_IWL<25149> A_IWL<25148> A_IWL<25147> A_IWL<25146> A_IWL<25145> A_IWL<25144> A_IWL<25143> A_IWL<25142> A_IWL<25141> A_IWL<25140> A_IWL<25139> A_IWL<25138> A_IWL<25137> A_IWL<25136> A_IWL<25135> A_IWL<25134> A_IWL<25133> A_IWL<25132> A_IWL<25131> A_IWL<25130> A_IWL<25129> A_IWL<25128> A_IWL<25127> A_IWL<25126> A_IWL<25125> A_IWL<25124> A_IWL<25123> A_IWL<25122> A_IWL<25121> A_IWL<25120> A_IWL<25119> A_IWL<25118> A_IWL<25117> A_IWL<25116> A_IWL<25115> A_IWL<25114> A_IWL<25113> A_IWL<25112> A_IWL<25111> A_IWL<25110> A_IWL<25109> A_IWL<25108> A_IWL<25107> A_IWL<25106> A_IWL<25105> A_IWL<25104> A_IWL<25103> A_IWL<25102> A_IWL<25101> A_IWL<25100> A_IWL<25099> A_IWL<25098> A_IWL<25097> A_IWL<25096> A_IWL<25095> A_IWL<25094> A_IWL<25093> A_IWL<25092> A_IWL<25091> A_IWL<25090> A_IWL<25089> A_IWL<25088> A_IWL<26111> A_IWL<26110> A_IWL<26109> A_IWL<26108> A_IWL<26107> A_IWL<26106> A_IWL<26105> A_IWL<26104> A_IWL<26103> A_IWL<26102> A_IWL<26101> A_IWL<26100> A_IWL<26099> A_IWL<26098> A_IWL<26097> A_IWL<26096> A_IWL<26095> A_IWL<26094> A_IWL<26093> A_IWL<26092> A_IWL<26091> A_IWL<26090> A_IWL<26089> A_IWL<26088> A_IWL<26087> A_IWL<26086> A_IWL<26085> A_IWL<26084> A_IWL<26083> A_IWL<26082> A_IWL<26081> A_IWL<26080> A_IWL<26079> A_IWL<26078> A_IWL<26077> A_IWL<26076> A_IWL<26075> A_IWL<26074> A_IWL<26073> A_IWL<26072> A_IWL<26071> A_IWL<26070> A_IWL<26069> A_IWL<26068> A_IWL<26067> A_IWL<26066> A_IWL<26065> A_IWL<26064> A_IWL<26063> A_IWL<26062> A_IWL<26061> A_IWL<26060> A_IWL<26059> A_IWL<26058> A_IWL<26057> A_IWL<26056> A_IWL<26055> A_IWL<26054> A_IWL<26053> A_IWL<26052> A_IWL<26051> A_IWL<26050> A_IWL<26049> A_IWL<26048> A_IWL<26047> A_IWL<26046> A_IWL<26045> A_IWL<26044> A_IWL<26043> A_IWL<26042> A_IWL<26041> A_IWL<26040> A_IWL<26039> A_IWL<26038> A_IWL<26037> A_IWL<26036> A_IWL<26035> A_IWL<26034> A_IWL<26033> A_IWL<26032> A_IWL<26031> A_IWL<26030> A_IWL<26029> A_IWL<26028> A_IWL<26027> A_IWL<26026> A_IWL<26025> A_IWL<26024> A_IWL<26023> A_IWL<26022> A_IWL<26021> A_IWL<26020> A_IWL<26019> A_IWL<26018> A_IWL<26017> A_IWL<26016> A_IWL<26015> A_IWL<26014> A_IWL<26013> A_IWL<26012> A_IWL<26011> A_IWL<26010> A_IWL<26009> A_IWL<26008> A_IWL<26007> A_IWL<26006> A_IWL<26005> A_IWL<26004> A_IWL<26003> A_IWL<26002> A_IWL<26001> A_IWL<26000> A_IWL<25999> A_IWL<25998> A_IWL<25997> A_IWL<25996> A_IWL<25995> A_IWL<25994> A_IWL<25993> A_IWL<25992> A_IWL<25991> A_IWL<25990> A_IWL<25989> A_IWL<25988> A_IWL<25987> A_IWL<25986> A_IWL<25985> A_IWL<25984> A_IWL<25983> A_IWL<25982> A_IWL<25981> A_IWL<25980> A_IWL<25979> A_IWL<25978> A_IWL<25977> A_IWL<25976> A_IWL<25975> A_IWL<25974> A_IWL<25973> A_IWL<25972> A_IWL<25971> A_IWL<25970> A_IWL<25969> A_IWL<25968> A_IWL<25967> A_IWL<25966> A_IWL<25965> A_IWL<25964> A_IWL<25963> A_IWL<25962> A_IWL<25961> A_IWL<25960> A_IWL<25959> A_IWL<25958> A_IWL<25957> A_IWL<25956> A_IWL<25955> A_IWL<25954> A_IWL<25953> A_IWL<25952> A_IWL<25951> A_IWL<25950> A_IWL<25949> A_IWL<25948> A_IWL<25947> A_IWL<25946> A_IWL<25945> A_IWL<25944> A_IWL<25943> A_IWL<25942> A_IWL<25941> A_IWL<25940> A_IWL<25939> A_IWL<25938> A_IWL<25937> A_IWL<25936> A_IWL<25935> A_IWL<25934> A_IWL<25933> A_IWL<25932> A_IWL<25931> A_IWL<25930> A_IWL<25929> A_IWL<25928> A_IWL<25927> A_IWL<25926> A_IWL<25925> A_IWL<25924> A_IWL<25923> A_IWL<25922> A_IWL<25921> A_IWL<25920> A_IWL<25919> A_IWL<25918> A_IWL<25917> A_IWL<25916> A_IWL<25915> A_IWL<25914> A_IWL<25913> A_IWL<25912> A_IWL<25911> A_IWL<25910> A_IWL<25909> A_IWL<25908> A_IWL<25907> A_IWL<25906> A_IWL<25905> A_IWL<25904> A_IWL<25903> A_IWL<25902> A_IWL<25901> A_IWL<25900> A_IWL<25899> A_IWL<25898> A_IWL<25897> A_IWL<25896> A_IWL<25895> A_IWL<25894> A_IWL<25893> A_IWL<25892> A_IWL<25891> A_IWL<25890> A_IWL<25889> A_IWL<25888> A_IWL<25887> A_IWL<25886> A_IWL<25885> A_IWL<25884> A_IWL<25883> A_IWL<25882> A_IWL<25881> A_IWL<25880> A_IWL<25879> A_IWL<25878> A_IWL<25877> A_IWL<25876> A_IWL<25875> A_IWL<25874> A_IWL<25873> A_IWL<25872> A_IWL<25871> A_IWL<25870> A_IWL<25869> A_IWL<25868> A_IWL<25867> A_IWL<25866> A_IWL<25865> A_IWL<25864> A_IWL<25863> A_IWL<25862> A_IWL<25861> A_IWL<25860> A_IWL<25859> A_IWL<25858> A_IWL<25857> A_IWL<25856> A_IWL<25855> A_IWL<25854> A_IWL<25853> A_IWL<25852> A_IWL<25851> A_IWL<25850> A_IWL<25849> A_IWL<25848> A_IWL<25847> A_IWL<25846> A_IWL<25845> A_IWL<25844> A_IWL<25843> A_IWL<25842> A_IWL<25841> A_IWL<25840> A_IWL<25839> A_IWL<25838> A_IWL<25837> A_IWL<25836> A_IWL<25835> A_IWL<25834> A_IWL<25833> A_IWL<25832> A_IWL<25831> A_IWL<25830> A_IWL<25829> A_IWL<25828> A_IWL<25827> A_IWL<25826> A_IWL<25825> A_IWL<25824> A_IWL<25823> A_IWL<25822> A_IWL<25821> A_IWL<25820> A_IWL<25819> A_IWL<25818> A_IWL<25817> A_IWL<25816> A_IWL<25815> A_IWL<25814> A_IWL<25813> A_IWL<25812> A_IWL<25811> A_IWL<25810> A_IWL<25809> A_IWL<25808> A_IWL<25807> A_IWL<25806> A_IWL<25805> A_IWL<25804> A_IWL<25803> A_IWL<25802> A_IWL<25801> A_IWL<25800> A_IWL<25799> A_IWL<25798> A_IWL<25797> A_IWL<25796> A_IWL<25795> A_IWL<25794> A_IWL<25793> A_IWL<25792> A_IWL<25791> A_IWL<25790> A_IWL<25789> A_IWL<25788> A_IWL<25787> A_IWL<25786> A_IWL<25785> A_IWL<25784> A_IWL<25783> A_IWL<25782> A_IWL<25781> A_IWL<25780> A_IWL<25779> A_IWL<25778> A_IWL<25777> A_IWL<25776> A_IWL<25775> A_IWL<25774> A_IWL<25773> A_IWL<25772> A_IWL<25771> A_IWL<25770> A_IWL<25769> A_IWL<25768> A_IWL<25767> A_IWL<25766> A_IWL<25765> A_IWL<25764> A_IWL<25763> A_IWL<25762> A_IWL<25761> A_IWL<25760> A_IWL<25759> A_IWL<25758> A_IWL<25757> A_IWL<25756> A_IWL<25755> A_IWL<25754> A_IWL<25753> A_IWL<25752> A_IWL<25751> A_IWL<25750> A_IWL<25749> A_IWL<25748> A_IWL<25747> A_IWL<25746> A_IWL<25745> A_IWL<25744> A_IWL<25743> A_IWL<25742> A_IWL<25741> A_IWL<25740> A_IWL<25739> A_IWL<25738> A_IWL<25737> A_IWL<25736> A_IWL<25735> A_IWL<25734> A_IWL<25733> A_IWL<25732> A_IWL<25731> A_IWL<25730> A_IWL<25729> A_IWL<25728> A_IWL<25727> A_IWL<25726> A_IWL<25725> A_IWL<25724> A_IWL<25723> A_IWL<25722> A_IWL<25721> A_IWL<25720> A_IWL<25719> A_IWL<25718> A_IWL<25717> A_IWL<25716> A_IWL<25715> A_IWL<25714> A_IWL<25713> A_IWL<25712> A_IWL<25711> A_IWL<25710> A_IWL<25709> A_IWL<25708> A_IWL<25707> A_IWL<25706> A_IWL<25705> A_IWL<25704> A_IWL<25703> A_IWL<25702> A_IWL<25701> A_IWL<25700> A_IWL<25699> A_IWL<25698> A_IWL<25697> A_IWL<25696> A_IWL<25695> A_IWL<25694> A_IWL<25693> A_IWL<25692> A_IWL<25691> A_IWL<25690> A_IWL<25689> A_IWL<25688> A_IWL<25687> A_IWL<25686> A_IWL<25685> A_IWL<25684> A_IWL<25683> A_IWL<25682> A_IWL<25681> A_IWL<25680> A_IWL<25679> A_IWL<25678> A_IWL<25677> A_IWL<25676> A_IWL<25675> A_IWL<25674> A_IWL<25673> A_IWL<25672> A_IWL<25671> A_IWL<25670> A_IWL<25669> A_IWL<25668> A_IWL<25667> A_IWL<25666> A_IWL<25665> A_IWL<25664> A_IWL<25663> A_IWL<25662> A_IWL<25661> A_IWL<25660> A_IWL<25659> A_IWL<25658> A_IWL<25657> A_IWL<25656> A_IWL<25655> A_IWL<25654> A_IWL<25653> A_IWL<25652> A_IWL<25651> A_IWL<25650> A_IWL<25649> A_IWL<25648> A_IWL<25647> A_IWL<25646> A_IWL<25645> A_IWL<25644> A_IWL<25643> A_IWL<25642> A_IWL<25641> A_IWL<25640> A_IWL<25639> A_IWL<25638> A_IWL<25637> A_IWL<25636> A_IWL<25635> A_IWL<25634> A_IWL<25633> A_IWL<25632> A_IWL<25631> A_IWL<25630> A_IWL<25629> A_IWL<25628> A_IWL<25627> A_IWL<25626> A_IWL<25625> A_IWL<25624> A_IWL<25623> A_IWL<25622> A_IWL<25621> A_IWL<25620> A_IWL<25619> A_IWL<25618> A_IWL<25617> A_IWL<25616> A_IWL<25615> A_IWL<25614> A_IWL<25613> A_IWL<25612> A_IWL<25611> A_IWL<25610> A_IWL<25609> A_IWL<25608> A_IWL<25607> A_IWL<25606> A_IWL<25605> A_IWL<25604> A_IWL<25603> A_IWL<25602> A_IWL<25601> A_IWL<25600> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<49> A_BLC<99> A_BLC<98> A_BLC_TOP<99> A_BLC_TOP<98> A_BLT<99> A_BLT<98> A_BLT_TOP<99> A_BLT_TOP<98> A_IWL<25087> A_IWL<25086> A_IWL<25085> A_IWL<25084> A_IWL<25083> A_IWL<25082> A_IWL<25081> A_IWL<25080> A_IWL<25079> A_IWL<25078> A_IWL<25077> A_IWL<25076> A_IWL<25075> A_IWL<25074> A_IWL<25073> A_IWL<25072> A_IWL<25071> A_IWL<25070> A_IWL<25069> A_IWL<25068> A_IWL<25067> A_IWL<25066> A_IWL<25065> A_IWL<25064> A_IWL<25063> A_IWL<25062> A_IWL<25061> A_IWL<25060> A_IWL<25059> A_IWL<25058> A_IWL<25057> A_IWL<25056> A_IWL<25055> A_IWL<25054> A_IWL<25053> A_IWL<25052> A_IWL<25051> A_IWL<25050> A_IWL<25049> A_IWL<25048> A_IWL<25047> A_IWL<25046> A_IWL<25045> A_IWL<25044> A_IWL<25043> A_IWL<25042> A_IWL<25041> A_IWL<25040> A_IWL<25039> A_IWL<25038> A_IWL<25037> A_IWL<25036> A_IWL<25035> A_IWL<25034> A_IWL<25033> A_IWL<25032> A_IWL<25031> A_IWL<25030> A_IWL<25029> A_IWL<25028> A_IWL<25027> A_IWL<25026> A_IWL<25025> A_IWL<25024> A_IWL<25023> A_IWL<25022> A_IWL<25021> A_IWL<25020> A_IWL<25019> A_IWL<25018> A_IWL<25017> A_IWL<25016> A_IWL<25015> A_IWL<25014> A_IWL<25013> A_IWL<25012> A_IWL<25011> A_IWL<25010> A_IWL<25009> A_IWL<25008> A_IWL<25007> A_IWL<25006> A_IWL<25005> A_IWL<25004> A_IWL<25003> A_IWL<25002> A_IWL<25001> A_IWL<25000> A_IWL<24999> A_IWL<24998> A_IWL<24997> A_IWL<24996> A_IWL<24995> A_IWL<24994> A_IWL<24993> A_IWL<24992> A_IWL<24991> A_IWL<24990> A_IWL<24989> A_IWL<24988> A_IWL<24987> A_IWL<24986> A_IWL<24985> A_IWL<24984> A_IWL<24983> A_IWL<24982> A_IWL<24981> A_IWL<24980> A_IWL<24979> A_IWL<24978> A_IWL<24977> A_IWL<24976> A_IWL<24975> A_IWL<24974> A_IWL<24973> A_IWL<24972> A_IWL<24971> A_IWL<24970> A_IWL<24969> A_IWL<24968> A_IWL<24967> A_IWL<24966> A_IWL<24965> A_IWL<24964> A_IWL<24963> A_IWL<24962> A_IWL<24961> A_IWL<24960> A_IWL<24959> A_IWL<24958> A_IWL<24957> A_IWL<24956> A_IWL<24955> A_IWL<24954> A_IWL<24953> A_IWL<24952> A_IWL<24951> A_IWL<24950> A_IWL<24949> A_IWL<24948> A_IWL<24947> A_IWL<24946> A_IWL<24945> A_IWL<24944> A_IWL<24943> A_IWL<24942> A_IWL<24941> A_IWL<24940> A_IWL<24939> A_IWL<24938> A_IWL<24937> A_IWL<24936> A_IWL<24935> A_IWL<24934> A_IWL<24933> A_IWL<24932> A_IWL<24931> A_IWL<24930> A_IWL<24929> A_IWL<24928> A_IWL<24927> A_IWL<24926> A_IWL<24925> A_IWL<24924> A_IWL<24923> A_IWL<24922> A_IWL<24921> A_IWL<24920> A_IWL<24919> A_IWL<24918> A_IWL<24917> A_IWL<24916> A_IWL<24915> A_IWL<24914> A_IWL<24913> A_IWL<24912> A_IWL<24911> A_IWL<24910> A_IWL<24909> A_IWL<24908> A_IWL<24907> A_IWL<24906> A_IWL<24905> A_IWL<24904> A_IWL<24903> A_IWL<24902> A_IWL<24901> A_IWL<24900> A_IWL<24899> A_IWL<24898> A_IWL<24897> A_IWL<24896> A_IWL<24895> A_IWL<24894> A_IWL<24893> A_IWL<24892> A_IWL<24891> A_IWL<24890> A_IWL<24889> A_IWL<24888> A_IWL<24887> A_IWL<24886> A_IWL<24885> A_IWL<24884> A_IWL<24883> A_IWL<24882> A_IWL<24881> A_IWL<24880> A_IWL<24879> A_IWL<24878> A_IWL<24877> A_IWL<24876> A_IWL<24875> A_IWL<24874> A_IWL<24873> A_IWL<24872> A_IWL<24871> A_IWL<24870> A_IWL<24869> A_IWL<24868> A_IWL<24867> A_IWL<24866> A_IWL<24865> A_IWL<24864> A_IWL<24863> A_IWL<24862> A_IWL<24861> A_IWL<24860> A_IWL<24859> A_IWL<24858> A_IWL<24857> A_IWL<24856> A_IWL<24855> A_IWL<24854> A_IWL<24853> A_IWL<24852> A_IWL<24851> A_IWL<24850> A_IWL<24849> A_IWL<24848> A_IWL<24847> A_IWL<24846> A_IWL<24845> A_IWL<24844> A_IWL<24843> A_IWL<24842> A_IWL<24841> A_IWL<24840> A_IWL<24839> A_IWL<24838> A_IWL<24837> A_IWL<24836> A_IWL<24835> A_IWL<24834> A_IWL<24833> A_IWL<24832> A_IWL<24831> A_IWL<24830> A_IWL<24829> A_IWL<24828> A_IWL<24827> A_IWL<24826> A_IWL<24825> A_IWL<24824> A_IWL<24823> A_IWL<24822> A_IWL<24821> A_IWL<24820> A_IWL<24819> A_IWL<24818> A_IWL<24817> A_IWL<24816> A_IWL<24815> A_IWL<24814> A_IWL<24813> A_IWL<24812> A_IWL<24811> A_IWL<24810> A_IWL<24809> A_IWL<24808> A_IWL<24807> A_IWL<24806> A_IWL<24805> A_IWL<24804> A_IWL<24803> A_IWL<24802> A_IWL<24801> A_IWL<24800> A_IWL<24799> A_IWL<24798> A_IWL<24797> A_IWL<24796> A_IWL<24795> A_IWL<24794> A_IWL<24793> A_IWL<24792> A_IWL<24791> A_IWL<24790> A_IWL<24789> A_IWL<24788> A_IWL<24787> A_IWL<24786> A_IWL<24785> A_IWL<24784> A_IWL<24783> A_IWL<24782> A_IWL<24781> A_IWL<24780> A_IWL<24779> A_IWL<24778> A_IWL<24777> A_IWL<24776> A_IWL<24775> A_IWL<24774> A_IWL<24773> A_IWL<24772> A_IWL<24771> A_IWL<24770> A_IWL<24769> A_IWL<24768> A_IWL<24767> A_IWL<24766> A_IWL<24765> A_IWL<24764> A_IWL<24763> A_IWL<24762> A_IWL<24761> A_IWL<24760> A_IWL<24759> A_IWL<24758> A_IWL<24757> A_IWL<24756> A_IWL<24755> A_IWL<24754> A_IWL<24753> A_IWL<24752> A_IWL<24751> A_IWL<24750> A_IWL<24749> A_IWL<24748> A_IWL<24747> A_IWL<24746> A_IWL<24745> A_IWL<24744> A_IWL<24743> A_IWL<24742> A_IWL<24741> A_IWL<24740> A_IWL<24739> A_IWL<24738> A_IWL<24737> A_IWL<24736> A_IWL<24735> A_IWL<24734> A_IWL<24733> A_IWL<24732> A_IWL<24731> A_IWL<24730> A_IWL<24729> A_IWL<24728> A_IWL<24727> A_IWL<24726> A_IWL<24725> A_IWL<24724> A_IWL<24723> A_IWL<24722> A_IWL<24721> A_IWL<24720> A_IWL<24719> A_IWL<24718> A_IWL<24717> A_IWL<24716> A_IWL<24715> A_IWL<24714> A_IWL<24713> A_IWL<24712> A_IWL<24711> A_IWL<24710> A_IWL<24709> A_IWL<24708> A_IWL<24707> A_IWL<24706> A_IWL<24705> A_IWL<24704> A_IWL<24703> A_IWL<24702> A_IWL<24701> A_IWL<24700> A_IWL<24699> A_IWL<24698> A_IWL<24697> A_IWL<24696> A_IWL<24695> A_IWL<24694> A_IWL<24693> A_IWL<24692> A_IWL<24691> A_IWL<24690> A_IWL<24689> A_IWL<24688> A_IWL<24687> A_IWL<24686> A_IWL<24685> A_IWL<24684> A_IWL<24683> A_IWL<24682> A_IWL<24681> A_IWL<24680> A_IWL<24679> A_IWL<24678> A_IWL<24677> A_IWL<24676> A_IWL<24675> A_IWL<24674> A_IWL<24673> A_IWL<24672> A_IWL<24671> A_IWL<24670> A_IWL<24669> A_IWL<24668> A_IWL<24667> A_IWL<24666> A_IWL<24665> A_IWL<24664> A_IWL<24663> A_IWL<24662> A_IWL<24661> A_IWL<24660> A_IWL<24659> A_IWL<24658> A_IWL<24657> A_IWL<24656> A_IWL<24655> A_IWL<24654> A_IWL<24653> A_IWL<24652> A_IWL<24651> A_IWL<24650> A_IWL<24649> A_IWL<24648> A_IWL<24647> A_IWL<24646> A_IWL<24645> A_IWL<24644> A_IWL<24643> A_IWL<24642> A_IWL<24641> A_IWL<24640> A_IWL<24639> A_IWL<24638> A_IWL<24637> A_IWL<24636> A_IWL<24635> A_IWL<24634> A_IWL<24633> A_IWL<24632> A_IWL<24631> A_IWL<24630> A_IWL<24629> A_IWL<24628> A_IWL<24627> A_IWL<24626> A_IWL<24625> A_IWL<24624> A_IWL<24623> A_IWL<24622> A_IWL<24621> A_IWL<24620> A_IWL<24619> A_IWL<24618> A_IWL<24617> A_IWL<24616> A_IWL<24615> A_IWL<24614> A_IWL<24613> A_IWL<24612> A_IWL<24611> A_IWL<24610> A_IWL<24609> A_IWL<24608> A_IWL<24607> A_IWL<24606> A_IWL<24605> A_IWL<24604> A_IWL<24603> A_IWL<24602> A_IWL<24601> A_IWL<24600> A_IWL<24599> A_IWL<24598> A_IWL<24597> A_IWL<24596> A_IWL<24595> A_IWL<24594> A_IWL<24593> A_IWL<24592> A_IWL<24591> A_IWL<24590> A_IWL<24589> A_IWL<24588> A_IWL<24587> A_IWL<24586> A_IWL<24585> A_IWL<24584> A_IWL<24583> A_IWL<24582> A_IWL<24581> A_IWL<24580> A_IWL<24579> A_IWL<24578> A_IWL<24577> A_IWL<24576> A_IWL<25599> A_IWL<25598> A_IWL<25597> A_IWL<25596> A_IWL<25595> A_IWL<25594> A_IWL<25593> A_IWL<25592> A_IWL<25591> A_IWL<25590> A_IWL<25589> A_IWL<25588> A_IWL<25587> A_IWL<25586> A_IWL<25585> A_IWL<25584> A_IWL<25583> A_IWL<25582> A_IWL<25581> A_IWL<25580> A_IWL<25579> A_IWL<25578> A_IWL<25577> A_IWL<25576> A_IWL<25575> A_IWL<25574> A_IWL<25573> A_IWL<25572> A_IWL<25571> A_IWL<25570> A_IWL<25569> A_IWL<25568> A_IWL<25567> A_IWL<25566> A_IWL<25565> A_IWL<25564> A_IWL<25563> A_IWL<25562> A_IWL<25561> A_IWL<25560> A_IWL<25559> A_IWL<25558> A_IWL<25557> A_IWL<25556> A_IWL<25555> A_IWL<25554> A_IWL<25553> A_IWL<25552> A_IWL<25551> A_IWL<25550> A_IWL<25549> A_IWL<25548> A_IWL<25547> A_IWL<25546> A_IWL<25545> A_IWL<25544> A_IWL<25543> A_IWL<25542> A_IWL<25541> A_IWL<25540> A_IWL<25539> A_IWL<25538> A_IWL<25537> A_IWL<25536> A_IWL<25535> A_IWL<25534> A_IWL<25533> A_IWL<25532> A_IWL<25531> A_IWL<25530> A_IWL<25529> A_IWL<25528> A_IWL<25527> A_IWL<25526> A_IWL<25525> A_IWL<25524> A_IWL<25523> A_IWL<25522> A_IWL<25521> A_IWL<25520> A_IWL<25519> A_IWL<25518> A_IWL<25517> A_IWL<25516> A_IWL<25515> A_IWL<25514> A_IWL<25513> A_IWL<25512> A_IWL<25511> A_IWL<25510> A_IWL<25509> A_IWL<25508> A_IWL<25507> A_IWL<25506> A_IWL<25505> A_IWL<25504> A_IWL<25503> A_IWL<25502> A_IWL<25501> A_IWL<25500> A_IWL<25499> A_IWL<25498> A_IWL<25497> A_IWL<25496> A_IWL<25495> A_IWL<25494> A_IWL<25493> A_IWL<25492> A_IWL<25491> A_IWL<25490> A_IWL<25489> A_IWL<25488> A_IWL<25487> A_IWL<25486> A_IWL<25485> A_IWL<25484> A_IWL<25483> A_IWL<25482> A_IWL<25481> A_IWL<25480> A_IWL<25479> A_IWL<25478> A_IWL<25477> A_IWL<25476> A_IWL<25475> A_IWL<25474> A_IWL<25473> A_IWL<25472> A_IWL<25471> A_IWL<25470> A_IWL<25469> A_IWL<25468> A_IWL<25467> A_IWL<25466> A_IWL<25465> A_IWL<25464> A_IWL<25463> A_IWL<25462> A_IWL<25461> A_IWL<25460> A_IWL<25459> A_IWL<25458> A_IWL<25457> A_IWL<25456> A_IWL<25455> A_IWL<25454> A_IWL<25453> A_IWL<25452> A_IWL<25451> A_IWL<25450> A_IWL<25449> A_IWL<25448> A_IWL<25447> A_IWL<25446> A_IWL<25445> A_IWL<25444> A_IWL<25443> A_IWL<25442> A_IWL<25441> A_IWL<25440> A_IWL<25439> A_IWL<25438> A_IWL<25437> A_IWL<25436> A_IWL<25435> A_IWL<25434> A_IWL<25433> A_IWL<25432> A_IWL<25431> A_IWL<25430> A_IWL<25429> A_IWL<25428> A_IWL<25427> A_IWL<25426> A_IWL<25425> A_IWL<25424> A_IWL<25423> A_IWL<25422> A_IWL<25421> A_IWL<25420> A_IWL<25419> A_IWL<25418> A_IWL<25417> A_IWL<25416> A_IWL<25415> A_IWL<25414> A_IWL<25413> A_IWL<25412> A_IWL<25411> A_IWL<25410> A_IWL<25409> A_IWL<25408> A_IWL<25407> A_IWL<25406> A_IWL<25405> A_IWL<25404> A_IWL<25403> A_IWL<25402> A_IWL<25401> A_IWL<25400> A_IWL<25399> A_IWL<25398> A_IWL<25397> A_IWL<25396> A_IWL<25395> A_IWL<25394> A_IWL<25393> A_IWL<25392> A_IWL<25391> A_IWL<25390> A_IWL<25389> A_IWL<25388> A_IWL<25387> A_IWL<25386> A_IWL<25385> A_IWL<25384> A_IWL<25383> A_IWL<25382> A_IWL<25381> A_IWL<25380> A_IWL<25379> A_IWL<25378> A_IWL<25377> A_IWL<25376> A_IWL<25375> A_IWL<25374> A_IWL<25373> A_IWL<25372> A_IWL<25371> A_IWL<25370> A_IWL<25369> A_IWL<25368> A_IWL<25367> A_IWL<25366> A_IWL<25365> A_IWL<25364> A_IWL<25363> A_IWL<25362> A_IWL<25361> A_IWL<25360> A_IWL<25359> A_IWL<25358> A_IWL<25357> A_IWL<25356> A_IWL<25355> A_IWL<25354> A_IWL<25353> A_IWL<25352> A_IWL<25351> A_IWL<25350> A_IWL<25349> A_IWL<25348> A_IWL<25347> A_IWL<25346> A_IWL<25345> A_IWL<25344> A_IWL<25343> A_IWL<25342> A_IWL<25341> A_IWL<25340> A_IWL<25339> A_IWL<25338> A_IWL<25337> A_IWL<25336> A_IWL<25335> A_IWL<25334> A_IWL<25333> A_IWL<25332> A_IWL<25331> A_IWL<25330> A_IWL<25329> A_IWL<25328> A_IWL<25327> A_IWL<25326> A_IWL<25325> A_IWL<25324> A_IWL<25323> A_IWL<25322> A_IWL<25321> A_IWL<25320> A_IWL<25319> A_IWL<25318> A_IWL<25317> A_IWL<25316> A_IWL<25315> A_IWL<25314> A_IWL<25313> A_IWL<25312> A_IWL<25311> A_IWL<25310> A_IWL<25309> A_IWL<25308> A_IWL<25307> A_IWL<25306> A_IWL<25305> A_IWL<25304> A_IWL<25303> A_IWL<25302> A_IWL<25301> A_IWL<25300> A_IWL<25299> A_IWL<25298> A_IWL<25297> A_IWL<25296> A_IWL<25295> A_IWL<25294> A_IWL<25293> A_IWL<25292> A_IWL<25291> A_IWL<25290> A_IWL<25289> A_IWL<25288> A_IWL<25287> A_IWL<25286> A_IWL<25285> A_IWL<25284> A_IWL<25283> A_IWL<25282> A_IWL<25281> A_IWL<25280> A_IWL<25279> A_IWL<25278> A_IWL<25277> A_IWL<25276> A_IWL<25275> A_IWL<25274> A_IWL<25273> A_IWL<25272> A_IWL<25271> A_IWL<25270> A_IWL<25269> A_IWL<25268> A_IWL<25267> A_IWL<25266> A_IWL<25265> A_IWL<25264> A_IWL<25263> A_IWL<25262> A_IWL<25261> A_IWL<25260> A_IWL<25259> A_IWL<25258> A_IWL<25257> A_IWL<25256> A_IWL<25255> A_IWL<25254> A_IWL<25253> A_IWL<25252> A_IWL<25251> A_IWL<25250> A_IWL<25249> A_IWL<25248> A_IWL<25247> A_IWL<25246> A_IWL<25245> A_IWL<25244> A_IWL<25243> A_IWL<25242> A_IWL<25241> A_IWL<25240> A_IWL<25239> A_IWL<25238> A_IWL<25237> A_IWL<25236> A_IWL<25235> A_IWL<25234> A_IWL<25233> A_IWL<25232> A_IWL<25231> A_IWL<25230> A_IWL<25229> A_IWL<25228> A_IWL<25227> A_IWL<25226> A_IWL<25225> A_IWL<25224> A_IWL<25223> A_IWL<25222> A_IWL<25221> A_IWL<25220> A_IWL<25219> A_IWL<25218> A_IWL<25217> A_IWL<25216> A_IWL<25215> A_IWL<25214> A_IWL<25213> A_IWL<25212> A_IWL<25211> A_IWL<25210> A_IWL<25209> A_IWL<25208> A_IWL<25207> A_IWL<25206> A_IWL<25205> A_IWL<25204> A_IWL<25203> A_IWL<25202> A_IWL<25201> A_IWL<25200> A_IWL<25199> A_IWL<25198> A_IWL<25197> A_IWL<25196> A_IWL<25195> A_IWL<25194> A_IWL<25193> A_IWL<25192> A_IWL<25191> A_IWL<25190> A_IWL<25189> A_IWL<25188> A_IWL<25187> A_IWL<25186> A_IWL<25185> A_IWL<25184> A_IWL<25183> A_IWL<25182> A_IWL<25181> A_IWL<25180> A_IWL<25179> A_IWL<25178> A_IWL<25177> A_IWL<25176> A_IWL<25175> A_IWL<25174> A_IWL<25173> A_IWL<25172> A_IWL<25171> A_IWL<25170> A_IWL<25169> A_IWL<25168> A_IWL<25167> A_IWL<25166> A_IWL<25165> A_IWL<25164> A_IWL<25163> A_IWL<25162> A_IWL<25161> A_IWL<25160> A_IWL<25159> A_IWL<25158> A_IWL<25157> A_IWL<25156> A_IWL<25155> A_IWL<25154> A_IWL<25153> A_IWL<25152> A_IWL<25151> A_IWL<25150> A_IWL<25149> A_IWL<25148> A_IWL<25147> A_IWL<25146> A_IWL<25145> A_IWL<25144> A_IWL<25143> A_IWL<25142> A_IWL<25141> A_IWL<25140> A_IWL<25139> A_IWL<25138> A_IWL<25137> A_IWL<25136> A_IWL<25135> A_IWL<25134> A_IWL<25133> A_IWL<25132> A_IWL<25131> A_IWL<25130> A_IWL<25129> A_IWL<25128> A_IWL<25127> A_IWL<25126> A_IWL<25125> A_IWL<25124> A_IWL<25123> A_IWL<25122> A_IWL<25121> A_IWL<25120> A_IWL<25119> A_IWL<25118> A_IWL<25117> A_IWL<25116> A_IWL<25115> A_IWL<25114> A_IWL<25113> A_IWL<25112> A_IWL<25111> A_IWL<25110> A_IWL<25109> A_IWL<25108> A_IWL<25107> A_IWL<25106> A_IWL<25105> A_IWL<25104> A_IWL<25103> A_IWL<25102> A_IWL<25101> A_IWL<25100> A_IWL<25099> A_IWL<25098> A_IWL<25097> A_IWL<25096> A_IWL<25095> A_IWL<25094> A_IWL<25093> A_IWL<25092> A_IWL<25091> A_IWL<25090> A_IWL<25089> A_IWL<25088> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<48> A_BLC<97> A_BLC<96> A_BLC_TOP<97> A_BLC_TOP<96> A_BLT<97> A_BLT<96> A_BLT_TOP<97> A_BLT_TOP<96> A_IWL<24575> A_IWL<24574> A_IWL<24573> A_IWL<24572> A_IWL<24571> A_IWL<24570> A_IWL<24569> A_IWL<24568> A_IWL<24567> A_IWL<24566> A_IWL<24565> A_IWL<24564> A_IWL<24563> A_IWL<24562> A_IWL<24561> A_IWL<24560> A_IWL<24559> A_IWL<24558> A_IWL<24557> A_IWL<24556> A_IWL<24555> A_IWL<24554> A_IWL<24553> A_IWL<24552> A_IWL<24551> A_IWL<24550> A_IWL<24549> A_IWL<24548> A_IWL<24547> A_IWL<24546> A_IWL<24545> A_IWL<24544> A_IWL<24543> A_IWL<24542> A_IWL<24541> A_IWL<24540> A_IWL<24539> A_IWL<24538> A_IWL<24537> A_IWL<24536> A_IWL<24535> A_IWL<24534> A_IWL<24533> A_IWL<24532> A_IWL<24531> A_IWL<24530> A_IWL<24529> A_IWL<24528> A_IWL<24527> A_IWL<24526> A_IWL<24525> A_IWL<24524> A_IWL<24523> A_IWL<24522> A_IWL<24521> A_IWL<24520> A_IWL<24519> A_IWL<24518> A_IWL<24517> A_IWL<24516> A_IWL<24515> A_IWL<24514> A_IWL<24513> A_IWL<24512> A_IWL<24511> A_IWL<24510> A_IWL<24509> A_IWL<24508> A_IWL<24507> A_IWL<24506> A_IWL<24505> A_IWL<24504> A_IWL<24503> A_IWL<24502> A_IWL<24501> A_IWL<24500> A_IWL<24499> A_IWL<24498> A_IWL<24497> A_IWL<24496> A_IWL<24495> A_IWL<24494> A_IWL<24493> A_IWL<24492> A_IWL<24491> A_IWL<24490> A_IWL<24489> A_IWL<24488> A_IWL<24487> A_IWL<24486> A_IWL<24485> A_IWL<24484> A_IWL<24483> A_IWL<24482> A_IWL<24481> A_IWL<24480> A_IWL<24479> A_IWL<24478> A_IWL<24477> A_IWL<24476> A_IWL<24475> A_IWL<24474> A_IWL<24473> A_IWL<24472> A_IWL<24471> A_IWL<24470> A_IWL<24469> A_IWL<24468> A_IWL<24467> A_IWL<24466> A_IWL<24465> A_IWL<24464> A_IWL<24463> A_IWL<24462> A_IWL<24461> A_IWL<24460> A_IWL<24459> A_IWL<24458> A_IWL<24457> A_IWL<24456> A_IWL<24455> A_IWL<24454> A_IWL<24453> A_IWL<24452> A_IWL<24451> A_IWL<24450> A_IWL<24449> A_IWL<24448> A_IWL<24447> A_IWL<24446> A_IWL<24445> A_IWL<24444> A_IWL<24443> A_IWL<24442> A_IWL<24441> A_IWL<24440> A_IWL<24439> A_IWL<24438> A_IWL<24437> A_IWL<24436> A_IWL<24435> A_IWL<24434> A_IWL<24433> A_IWL<24432> A_IWL<24431> A_IWL<24430> A_IWL<24429> A_IWL<24428> A_IWL<24427> A_IWL<24426> A_IWL<24425> A_IWL<24424> A_IWL<24423> A_IWL<24422> A_IWL<24421> A_IWL<24420> A_IWL<24419> A_IWL<24418> A_IWL<24417> A_IWL<24416> A_IWL<24415> A_IWL<24414> A_IWL<24413> A_IWL<24412> A_IWL<24411> A_IWL<24410> A_IWL<24409> A_IWL<24408> A_IWL<24407> A_IWL<24406> A_IWL<24405> A_IWL<24404> A_IWL<24403> A_IWL<24402> A_IWL<24401> A_IWL<24400> A_IWL<24399> A_IWL<24398> A_IWL<24397> A_IWL<24396> A_IWL<24395> A_IWL<24394> A_IWL<24393> A_IWL<24392> A_IWL<24391> A_IWL<24390> A_IWL<24389> A_IWL<24388> A_IWL<24387> A_IWL<24386> A_IWL<24385> A_IWL<24384> A_IWL<24383> A_IWL<24382> A_IWL<24381> A_IWL<24380> A_IWL<24379> A_IWL<24378> A_IWL<24377> A_IWL<24376> A_IWL<24375> A_IWL<24374> A_IWL<24373> A_IWL<24372> A_IWL<24371> A_IWL<24370> A_IWL<24369> A_IWL<24368> A_IWL<24367> A_IWL<24366> A_IWL<24365> A_IWL<24364> A_IWL<24363> A_IWL<24362> A_IWL<24361> A_IWL<24360> A_IWL<24359> A_IWL<24358> A_IWL<24357> A_IWL<24356> A_IWL<24355> A_IWL<24354> A_IWL<24353> A_IWL<24352> A_IWL<24351> A_IWL<24350> A_IWL<24349> A_IWL<24348> A_IWL<24347> A_IWL<24346> A_IWL<24345> A_IWL<24344> A_IWL<24343> A_IWL<24342> A_IWL<24341> A_IWL<24340> A_IWL<24339> A_IWL<24338> A_IWL<24337> A_IWL<24336> A_IWL<24335> A_IWL<24334> A_IWL<24333> A_IWL<24332> A_IWL<24331> A_IWL<24330> A_IWL<24329> A_IWL<24328> A_IWL<24327> A_IWL<24326> A_IWL<24325> A_IWL<24324> A_IWL<24323> A_IWL<24322> A_IWL<24321> A_IWL<24320> A_IWL<24319> A_IWL<24318> A_IWL<24317> A_IWL<24316> A_IWL<24315> A_IWL<24314> A_IWL<24313> A_IWL<24312> A_IWL<24311> A_IWL<24310> A_IWL<24309> A_IWL<24308> A_IWL<24307> A_IWL<24306> A_IWL<24305> A_IWL<24304> A_IWL<24303> A_IWL<24302> A_IWL<24301> A_IWL<24300> A_IWL<24299> A_IWL<24298> A_IWL<24297> A_IWL<24296> A_IWL<24295> A_IWL<24294> A_IWL<24293> A_IWL<24292> A_IWL<24291> A_IWL<24290> A_IWL<24289> A_IWL<24288> A_IWL<24287> A_IWL<24286> A_IWL<24285> A_IWL<24284> A_IWL<24283> A_IWL<24282> A_IWL<24281> A_IWL<24280> A_IWL<24279> A_IWL<24278> A_IWL<24277> A_IWL<24276> A_IWL<24275> A_IWL<24274> A_IWL<24273> A_IWL<24272> A_IWL<24271> A_IWL<24270> A_IWL<24269> A_IWL<24268> A_IWL<24267> A_IWL<24266> A_IWL<24265> A_IWL<24264> A_IWL<24263> A_IWL<24262> A_IWL<24261> A_IWL<24260> A_IWL<24259> A_IWL<24258> A_IWL<24257> A_IWL<24256> A_IWL<24255> A_IWL<24254> A_IWL<24253> A_IWL<24252> A_IWL<24251> A_IWL<24250> A_IWL<24249> A_IWL<24248> A_IWL<24247> A_IWL<24246> A_IWL<24245> A_IWL<24244> A_IWL<24243> A_IWL<24242> A_IWL<24241> A_IWL<24240> A_IWL<24239> A_IWL<24238> A_IWL<24237> A_IWL<24236> A_IWL<24235> A_IWL<24234> A_IWL<24233> A_IWL<24232> A_IWL<24231> A_IWL<24230> A_IWL<24229> A_IWL<24228> A_IWL<24227> A_IWL<24226> A_IWL<24225> A_IWL<24224> A_IWL<24223> A_IWL<24222> A_IWL<24221> A_IWL<24220> A_IWL<24219> A_IWL<24218> A_IWL<24217> A_IWL<24216> A_IWL<24215> A_IWL<24214> A_IWL<24213> A_IWL<24212> A_IWL<24211> A_IWL<24210> A_IWL<24209> A_IWL<24208> A_IWL<24207> A_IWL<24206> A_IWL<24205> A_IWL<24204> A_IWL<24203> A_IWL<24202> A_IWL<24201> A_IWL<24200> A_IWL<24199> A_IWL<24198> A_IWL<24197> A_IWL<24196> A_IWL<24195> A_IWL<24194> A_IWL<24193> A_IWL<24192> A_IWL<24191> A_IWL<24190> A_IWL<24189> A_IWL<24188> A_IWL<24187> A_IWL<24186> A_IWL<24185> A_IWL<24184> A_IWL<24183> A_IWL<24182> A_IWL<24181> A_IWL<24180> A_IWL<24179> A_IWL<24178> A_IWL<24177> A_IWL<24176> A_IWL<24175> A_IWL<24174> A_IWL<24173> A_IWL<24172> A_IWL<24171> A_IWL<24170> A_IWL<24169> A_IWL<24168> A_IWL<24167> A_IWL<24166> A_IWL<24165> A_IWL<24164> A_IWL<24163> A_IWL<24162> A_IWL<24161> A_IWL<24160> A_IWL<24159> A_IWL<24158> A_IWL<24157> A_IWL<24156> A_IWL<24155> A_IWL<24154> A_IWL<24153> A_IWL<24152> A_IWL<24151> A_IWL<24150> A_IWL<24149> A_IWL<24148> A_IWL<24147> A_IWL<24146> A_IWL<24145> A_IWL<24144> A_IWL<24143> A_IWL<24142> A_IWL<24141> A_IWL<24140> A_IWL<24139> A_IWL<24138> A_IWL<24137> A_IWL<24136> A_IWL<24135> A_IWL<24134> A_IWL<24133> A_IWL<24132> A_IWL<24131> A_IWL<24130> A_IWL<24129> A_IWL<24128> A_IWL<24127> A_IWL<24126> A_IWL<24125> A_IWL<24124> A_IWL<24123> A_IWL<24122> A_IWL<24121> A_IWL<24120> A_IWL<24119> A_IWL<24118> A_IWL<24117> A_IWL<24116> A_IWL<24115> A_IWL<24114> A_IWL<24113> A_IWL<24112> A_IWL<24111> A_IWL<24110> A_IWL<24109> A_IWL<24108> A_IWL<24107> A_IWL<24106> A_IWL<24105> A_IWL<24104> A_IWL<24103> A_IWL<24102> A_IWL<24101> A_IWL<24100> A_IWL<24099> A_IWL<24098> A_IWL<24097> A_IWL<24096> A_IWL<24095> A_IWL<24094> A_IWL<24093> A_IWL<24092> A_IWL<24091> A_IWL<24090> A_IWL<24089> A_IWL<24088> A_IWL<24087> A_IWL<24086> A_IWL<24085> A_IWL<24084> A_IWL<24083> A_IWL<24082> A_IWL<24081> A_IWL<24080> A_IWL<24079> A_IWL<24078> A_IWL<24077> A_IWL<24076> A_IWL<24075> A_IWL<24074> A_IWL<24073> A_IWL<24072> A_IWL<24071> A_IWL<24070> A_IWL<24069> A_IWL<24068> A_IWL<24067> A_IWL<24066> A_IWL<24065> A_IWL<24064> A_IWL<25087> A_IWL<25086> A_IWL<25085> A_IWL<25084> A_IWL<25083> A_IWL<25082> A_IWL<25081> A_IWL<25080> A_IWL<25079> A_IWL<25078> A_IWL<25077> A_IWL<25076> A_IWL<25075> A_IWL<25074> A_IWL<25073> A_IWL<25072> A_IWL<25071> A_IWL<25070> A_IWL<25069> A_IWL<25068> A_IWL<25067> A_IWL<25066> A_IWL<25065> A_IWL<25064> A_IWL<25063> A_IWL<25062> A_IWL<25061> A_IWL<25060> A_IWL<25059> A_IWL<25058> A_IWL<25057> A_IWL<25056> A_IWL<25055> A_IWL<25054> A_IWL<25053> A_IWL<25052> A_IWL<25051> A_IWL<25050> A_IWL<25049> A_IWL<25048> A_IWL<25047> A_IWL<25046> A_IWL<25045> A_IWL<25044> A_IWL<25043> A_IWL<25042> A_IWL<25041> A_IWL<25040> A_IWL<25039> A_IWL<25038> A_IWL<25037> A_IWL<25036> A_IWL<25035> A_IWL<25034> A_IWL<25033> A_IWL<25032> A_IWL<25031> A_IWL<25030> A_IWL<25029> A_IWL<25028> A_IWL<25027> A_IWL<25026> A_IWL<25025> A_IWL<25024> A_IWL<25023> A_IWL<25022> A_IWL<25021> A_IWL<25020> A_IWL<25019> A_IWL<25018> A_IWL<25017> A_IWL<25016> A_IWL<25015> A_IWL<25014> A_IWL<25013> A_IWL<25012> A_IWL<25011> A_IWL<25010> A_IWL<25009> A_IWL<25008> A_IWL<25007> A_IWL<25006> A_IWL<25005> A_IWL<25004> A_IWL<25003> A_IWL<25002> A_IWL<25001> A_IWL<25000> A_IWL<24999> A_IWL<24998> A_IWL<24997> A_IWL<24996> A_IWL<24995> A_IWL<24994> A_IWL<24993> A_IWL<24992> A_IWL<24991> A_IWL<24990> A_IWL<24989> A_IWL<24988> A_IWL<24987> A_IWL<24986> A_IWL<24985> A_IWL<24984> A_IWL<24983> A_IWL<24982> A_IWL<24981> A_IWL<24980> A_IWL<24979> A_IWL<24978> A_IWL<24977> A_IWL<24976> A_IWL<24975> A_IWL<24974> A_IWL<24973> A_IWL<24972> A_IWL<24971> A_IWL<24970> A_IWL<24969> A_IWL<24968> A_IWL<24967> A_IWL<24966> A_IWL<24965> A_IWL<24964> A_IWL<24963> A_IWL<24962> A_IWL<24961> A_IWL<24960> A_IWL<24959> A_IWL<24958> A_IWL<24957> A_IWL<24956> A_IWL<24955> A_IWL<24954> A_IWL<24953> A_IWL<24952> A_IWL<24951> A_IWL<24950> A_IWL<24949> A_IWL<24948> A_IWL<24947> A_IWL<24946> A_IWL<24945> A_IWL<24944> A_IWL<24943> A_IWL<24942> A_IWL<24941> A_IWL<24940> A_IWL<24939> A_IWL<24938> A_IWL<24937> A_IWL<24936> A_IWL<24935> A_IWL<24934> A_IWL<24933> A_IWL<24932> A_IWL<24931> A_IWL<24930> A_IWL<24929> A_IWL<24928> A_IWL<24927> A_IWL<24926> A_IWL<24925> A_IWL<24924> A_IWL<24923> A_IWL<24922> A_IWL<24921> A_IWL<24920> A_IWL<24919> A_IWL<24918> A_IWL<24917> A_IWL<24916> A_IWL<24915> A_IWL<24914> A_IWL<24913> A_IWL<24912> A_IWL<24911> A_IWL<24910> A_IWL<24909> A_IWL<24908> A_IWL<24907> A_IWL<24906> A_IWL<24905> A_IWL<24904> A_IWL<24903> A_IWL<24902> A_IWL<24901> A_IWL<24900> A_IWL<24899> A_IWL<24898> A_IWL<24897> A_IWL<24896> A_IWL<24895> A_IWL<24894> A_IWL<24893> A_IWL<24892> A_IWL<24891> A_IWL<24890> A_IWL<24889> A_IWL<24888> A_IWL<24887> A_IWL<24886> A_IWL<24885> A_IWL<24884> A_IWL<24883> A_IWL<24882> A_IWL<24881> A_IWL<24880> A_IWL<24879> A_IWL<24878> A_IWL<24877> A_IWL<24876> A_IWL<24875> A_IWL<24874> A_IWL<24873> A_IWL<24872> A_IWL<24871> A_IWL<24870> A_IWL<24869> A_IWL<24868> A_IWL<24867> A_IWL<24866> A_IWL<24865> A_IWL<24864> A_IWL<24863> A_IWL<24862> A_IWL<24861> A_IWL<24860> A_IWL<24859> A_IWL<24858> A_IWL<24857> A_IWL<24856> A_IWL<24855> A_IWL<24854> A_IWL<24853> A_IWL<24852> A_IWL<24851> A_IWL<24850> A_IWL<24849> A_IWL<24848> A_IWL<24847> A_IWL<24846> A_IWL<24845> A_IWL<24844> A_IWL<24843> A_IWL<24842> A_IWL<24841> A_IWL<24840> A_IWL<24839> A_IWL<24838> A_IWL<24837> A_IWL<24836> A_IWL<24835> A_IWL<24834> A_IWL<24833> A_IWL<24832> A_IWL<24831> A_IWL<24830> A_IWL<24829> A_IWL<24828> A_IWL<24827> A_IWL<24826> A_IWL<24825> A_IWL<24824> A_IWL<24823> A_IWL<24822> A_IWL<24821> A_IWL<24820> A_IWL<24819> A_IWL<24818> A_IWL<24817> A_IWL<24816> A_IWL<24815> A_IWL<24814> A_IWL<24813> A_IWL<24812> A_IWL<24811> A_IWL<24810> A_IWL<24809> A_IWL<24808> A_IWL<24807> A_IWL<24806> A_IWL<24805> A_IWL<24804> A_IWL<24803> A_IWL<24802> A_IWL<24801> A_IWL<24800> A_IWL<24799> A_IWL<24798> A_IWL<24797> A_IWL<24796> A_IWL<24795> A_IWL<24794> A_IWL<24793> A_IWL<24792> A_IWL<24791> A_IWL<24790> A_IWL<24789> A_IWL<24788> A_IWL<24787> A_IWL<24786> A_IWL<24785> A_IWL<24784> A_IWL<24783> A_IWL<24782> A_IWL<24781> A_IWL<24780> A_IWL<24779> A_IWL<24778> A_IWL<24777> A_IWL<24776> A_IWL<24775> A_IWL<24774> A_IWL<24773> A_IWL<24772> A_IWL<24771> A_IWL<24770> A_IWL<24769> A_IWL<24768> A_IWL<24767> A_IWL<24766> A_IWL<24765> A_IWL<24764> A_IWL<24763> A_IWL<24762> A_IWL<24761> A_IWL<24760> A_IWL<24759> A_IWL<24758> A_IWL<24757> A_IWL<24756> A_IWL<24755> A_IWL<24754> A_IWL<24753> A_IWL<24752> A_IWL<24751> A_IWL<24750> A_IWL<24749> A_IWL<24748> A_IWL<24747> A_IWL<24746> A_IWL<24745> A_IWL<24744> A_IWL<24743> A_IWL<24742> A_IWL<24741> A_IWL<24740> A_IWL<24739> A_IWL<24738> A_IWL<24737> A_IWL<24736> A_IWL<24735> A_IWL<24734> A_IWL<24733> A_IWL<24732> A_IWL<24731> A_IWL<24730> A_IWL<24729> A_IWL<24728> A_IWL<24727> A_IWL<24726> A_IWL<24725> A_IWL<24724> A_IWL<24723> A_IWL<24722> A_IWL<24721> A_IWL<24720> A_IWL<24719> A_IWL<24718> A_IWL<24717> A_IWL<24716> A_IWL<24715> A_IWL<24714> A_IWL<24713> A_IWL<24712> A_IWL<24711> A_IWL<24710> A_IWL<24709> A_IWL<24708> A_IWL<24707> A_IWL<24706> A_IWL<24705> A_IWL<24704> A_IWL<24703> A_IWL<24702> A_IWL<24701> A_IWL<24700> A_IWL<24699> A_IWL<24698> A_IWL<24697> A_IWL<24696> A_IWL<24695> A_IWL<24694> A_IWL<24693> A_IWL<24692> A_IWL<24691> A_IWL<24690> A_IWL<24689> A_IWL<24688> A_IWL<24687> A_IWL<24686> A_IWL<24685> A_IWL<24684> A_IWL<24683> A_IWL<24682> A_IWL<24681> A_IWL<24680> A_IWL<24679> A_IWL<24678> A_IWL<24677> A_IWL<24676> A_IWL<24675> A_IWL<24674> A_IWL<24673> A_IWL<24672> A_IWL<24671> A_IWL<24670> A_IWL<24669> A_IWL<24668> A_IWL<24667> A_IWL<24666> A_IWL<24665> A_IWL<24664> A_IWL<24663> A_IWL<24662> A_IWL<24661> A_IWL<24660> A_IWL<24659> A_IWL<24658> A_IWL<24657> A_IWL<24656> A_IWL<24655> A_IWL<24654> A_IWL<24653> A_IWL<24652> A_IWL<24651> A_IWL<24650> A_IWL<24649> A_IWL<24648> A_IWL<24647> A_IWL<24646> A_IWL<24645> A_IWL<24644> A_IWL<24643> A_IWL<24642> A_IWL<24641> A_IWL<24640> A_IWL<24639> A_IWL<24638> A_IWL<24637> A_IWL<24636> A_IWL<24635> A_IWL<24634> A_IWL<24633> A_IWL<24632> A_IWL<24631> A_IWL<24630> A_IWL<24629> A_IWL<24628> A_IWL<24627> A_IWL<24626> A_IWL<24625> A_IWL<24624> A_IWL<24623> A_IWL<24622> A_IWL<24621> A_IWL<24620> A_IWL<24619> A_IWL<24618> A_IWL<24617> A_IWL<24616> A_IWL<24615> A_IWL<24614> A_IWL<24613> A_IWL<24612> A_IWL<24611> A_IWL<24610> A_IWL<24609> A_IWL<24608> A_IWL<24607> A_IWL<24606> A_IWL<24605> A_IWL<24604> A_IWL<24603> A_IWL<24602> A_IWL<24601> A_IWL<24600> A_IWL<24599> A_IWL<24598> A_IWL<24597> A_IWL<24596> A_IWL<24595> A_IWL<24594> A_IWL<24593> A_IWL<24592> A_IWL<24591> A_IWL<24590> A_IWL<24589> A_IWL<24588> A_IWL<24587> A_IWL<24586> A_IWL<24585> A_IWL<24584> A_IWL<24583> A_IWL<24582> A_IWL<24581> A_IWL<24580> A_IWL<24579> A_IWL<24578> A_IWL<24577> A_IWL<24576> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<47> A_BLC<95> A_BLC<94> A_BLC_TOP<95> A_BLC_TOP<94> A_BLT<95> A_BLT<94> A_BLT_TOP<95> A_BLT_TOP<94> A_IWL<24063> A_IWL<24062> A_IWL<24061> A_IWL<24060> A_IWL<24059> A_IWL<24058> A_IWL<24057> A_IWL<24056> A_IWL<24055> A_IWL<24054> A_IWL<24053> A_IWL<24052> A_IWL<24051> A_IWL<24050> A_IWL<24049> A_IWL<24048> A_IWL<24047> A_IWL<24046> A_IWL<24045> A_IWL<24044> A_IWL<24043> A_IWL<24042> A_IWL<24041> A_IWL<24040> A_IWL<24039> A_IWL<24038> A_IWL<24037> A_IWL<24036> A_IWL<24035> A_IWL<24034> A_IWL<24033> A_IWL<24032> A_IWL<24031> A_IWL<24030> A_IWL<24029> A_IWL<24028> A_IWL<24027> A_IWL<24026> A_IWL<24025> A_IWL<24024> A_IWL<24023> A_IWL<24022> A_IWL<24021> A_IWL<24020> A_IWL<24019> A_IWL<24018> A_IWL<24017> A_IWL<24016> A_IWL<24015> A_IWL<24014> A_IWL<24013> A_IWL<24012> A_IWL<24011> A_IWL<24010> A_IWL<24009> A_IWL<24008> A_IWL<24007> A_IWL<24006> A_IWL<24005> A_IWL<24004> A_IWL<24003> A_IWL<24002> A_IWL<24001> A_IWL<24000> A_IWL<23999> A_IWL<23998> A_IWL<23997> A_IWL<23996> A_IWL<23995> A_IWL<23994> A_IWL<23993> A_IWL<23992> A_IWL<23991> A_IWL<23990> A_IWL<23989> A_IWL<23988> A_IWL<23987> A_IWL<23986> A_IWL<23985> A_IWL<23984> A_IWL<23983> A_IWL<23982> A_IWL<23981> A_IWL<23980> A_IWL<23979> A_IWL<23978> A_IWL<23977> A_IWL<23976> A_IWL<23975> A_IWL<23974> A_IWL<23973> A_IWL<23972> A_IWL<23971> A_IWL<23970> A_IWL<23969> A_IWL<23968> A_IWL<23967> A_IWL<23966> A_IWL<23965> A_IWL<23964> A_IWL<23963> A_IWL<23962> A_IWL<23961> A_IWL<23960> A_IWL<23959> A_IWL<23958> A_IWL<23957> A_IWL<23956> A_IWL<23955> A_IWL<23954> A_IWL<23953> A_IWL<23952> A_IWL<23951> A_IWL<23950> A_IWL<23949> A_IWL<23948> A_IWL<23947> A_IWL<23946> A_IWL<23945> A_IWL<23944> A_IWL<23943> A_IWL<23942> A_IWL<23941> A_IWL<23940> A_IWL<23939> A_IWL<23938> A_IWL<23937> A_IWL<23936> A_IWL<23935> A_IWL<23934> A_IWL<23933> A_IWL<23932> A_IWL<23931> A_IWL<23930> A_IWL<23929> A_IWL<23928> A_IWL<23927> A_IWL<23926> A_IWL<23925> A_IWL<23924> A_IWL<23923> A_IWL<23922> A_IWL<23921> A_IWL<23920> A_IWL<23919> A_IWL<23918> A_IWL<23917> A_IWL<23916> A_IWL<23915> A_IWL<23914> A_IWL<23913> A_IWL<23912> A_IWL<23911> A_IWL<23910> A_IWL<23909> A_IWL<23908> A_IWL<23907> A_IWL<23906> A_IWL<23905> A_IWL<23904> A_IWL<23903> A_IWL<23902> A_IWL<23901> A_IWL<23900> A_IWL<23899> A_IWL<23898> A_IWL<23897> A_IWL<23896> A_IWL<23895> A_IWL<23894> A_IWL<23893> A_IWL<23892> A_IWL<23891> A_IWL<23890> A_IWL<23889> A_IWL<23888> A_IWL<23887> A_IWL<23886> A_IWL<23885> A_IWL<23884> A_IWL<23883> A_IWL<23882> A_IWL<23881> A_IWL<23880> A_IWL<23879> A_IWL<23878> A_IWL<23877> A_IWL<23876> A_IWL<23875> A_IWL<23874> A_IWL<23873> A_IWL<23872> A_IWL<23871> A_IWL<23870> A_IWL<23869> A_IWL<23868> A_IWL<23867> A_IWL<23866> A_IWL<23865> A_IWL<23864> A_IWL<23863> A_IWL<23862> A_IWL<23861> A_IWL<23860> A_IWL<23859> A_IWL<23858> A_IWL<23857> A_IWL<23856> A_IWL<23855> A_IWL<23854> A_IWL<23853> A_IWL<23852> A_IWL<23851> A_IWL<23850> A_IWL<23849> A_IWL<23848> A_IWL<23847> A_IWL<23846> A_IWL<23845> A_IWL<23844> A_IWL<23843> A_IWL<23842> A_IWL<23841> A_IWL<23840> A_IWL<23839> A_IWL<23838> A_IWL<23837> A_IWL<23836> A_IWL<23835> A_IWL<23834> A_IWL<23833> A_IWL<23832> A_IWL<23831> A_IWL<23830> A_IWL<23829> A_IWL<23828> A_IWL<23827> A_IWL<23826> A_IWL<23825> A_IWL<23824> A_IWL<23823> A_IWL<23822> A_IWL<23821> A_IWL<23820> A_IWL<23819> A_IWL<23818> A_IWL<23817> A_IWL<23816> A_IWL<23815> A_IWL<23814> A_IWL<23813> A_IWL<23812> A_IWL<23811> A_IWL<23810> A_IWL<23809> A_IWL<23808> A_IWL<23807> A_IWL<23806> A_IWL<23805> A_IWL<23804> A_IWL<23803> A_IWL<23802> A_IWL<23801> A_IWL<23800> A_IWL<23799> A_IWL<23798> A_IWL<23797> A_IWL<23796> A_IWL<23795> A_IWL<23794> A_IWL<23793> A_IWL<23792> A_IWL<23791> A_IWL<23790> A_IWL<23789> A_IWL<23788> A_IWL<23787> A_IWL<23786> A_IWL<23785> A_IWL<23784> A_IWL<23783> A_IWL<23782> A_IWL<23781> A_IWL<23780> A_IWL<23779> A_IWL<23778> A_IWL<23777> A_IWL<23776> A_IWL<23775> A_IWL<23774> A_IWL<23773> A_IWL<23772> A_IWL<23771> A_IWL<23770> A_IWL<23769> A_IWL<23768> A_IWL<23767> A_IWL<23766> A_IWL<23765> A_IWL<23764> A_IWL<23763> A_IWL<23762> A_IWL<23761> A_IWL<23760> A_IWL<23759> A_IWL<23758> A_IWL<23757> A_IWL<23756> A_IWL<23755> A_IWL<23754> A_IWL<23753> A_IWL<23752> A_IWL<23751> A_IWL<23750> A_IWL<23749> A_IWL<23748> A_IWL<23747> A_IWL<23746> A_IWL<23745> A_IWL<23744> A_IWL<23743> A_IWL<23742> A_IWL<23741> A_IWL<23740> A_IWL<23739> A_IWL<23738> A_IWL<23737> A_IWL<23736> A_IWL<23735> A_IWL<23734> A_IWL<23733> A_IWL<23732> A_IWL<23731> A_IWL<23730> A_IWL<23729> A_IWL<23728> A_IWL<23727> A_IWL<23726> A_IWL<23725> A_IWL<23724> A_IWL<23723> A_IWL<23722> A_IWL<23721> A_IWL<23720> A_IWL<23719> A_IWL<23718> A_IWL<23717> A_IWL<23716> A_IWL<23715> A_IWL<23714> A_IWL<23713> A_IWL<23712> A_IWL<23711> A_IWL<23710> A_IWL<23709> A_IWL<23708> A_IWL<23707> A_IWL<23706> A_IWL<23705> A_IWL<23704> A_IWL<23703> A_IWL<23702> A_IWL<23701> A_IWL<23700> A_IWL<23699> A_IWL<23698> A_IWL<23697> A_IWL<23696> A_IWL<23695> A_IWL<23694> A_IWL<23693> A_IWL<23692> A_IWL<23691> A_IWL<23690> A_IWL<23689> A_IWL<23688> A_IWL<23687> A_IWL<23686> A_IWL<23685> A_IWL<23684> A_IWL<23683> A_IWL<23682> A_IWL<23681> A_IWL<23680> A_IWL<23679> A_IWL<23678> A_IWL<23677> A_IWL<23676> A_IWL<23675> A_IWL<23674> A_IWL<23673> A_IWL<23672> A_IWL<23671> A_IWL<23670> A_IWL<23669> A_IWL<23668> A_IWL<23667> A_IWL<23666> A_IWL<23665> A_IWL<23664> A_IWL<23663> A_IWL<23662> A_IWL<23661> A_IWL<23660> A_IWL<23659> A_IWL<23658> A_IWL<23657> A_IWL<23656> A_IWL<23655> A_IWL<23654> A_IWL<23653> A_IWL<23652> A_IWL<23651> A_IWL<23650> A_IWL<23649> A_IWL<23648> A_IWL<23647> A_IWL<23646> A_IWL<23645> A_IWL<23644> A_IWL<23643> A_IWL<23642> A_IWL<23641> A_IWL<23640> A_IWL<23639> A_IWL<23638> A_IWL<23637> A_IWL<23636> A_IWL<23635> A_IWL<23634> A_IWL<23633> A_IWL<23632> A_IWL<23631> A_IWL<23630> A_IWL<23629> A_IWL<23628> A_IWL<23627> A_IWL<23626> A_IWL<23625> A_IWL<23624> A_IWL<23623> A_IWL<23622> A_IWL<23621> A_IWL<23620> A_IWL<23619> A_IWL<23618> A_IWL<23617> A_IWL<23616> A_IWL<23615> A_IWL<23614> A_IWL<23613> A_IWL<23612> A_IWL<23611> A_IWL<23610> A_IWL<23609> A_IWL<23608> A_IWL<23607> A_IWL<23606> A_IWL<23605> A_IWL<23604> A_IWL<23603> A_IWL<23602> A_IWL<23601> A_IWL<23600> A_IWL<23599> A_IWL<23598> A_IWL<23597> A_IWL<23596> A_IWL<23595> A_IWL<23594> A_IWL<23593> A_IWL<23592> A_IWL<23591> A_IWL<23590> A_IWL<23589> A_IWL<23588> A_IWL<23587> A_IWL<23586> A_IWL<23585> A_IWL<23584> A_IWL<23583> A_IWL<23582> A_IWL<23581> A_IWL<23580> A_IWL<23579> A_IWL<23578> A_IWL<23577> A_IWL<23576> A_IWL<23575> A_IWL<23574> A_IWL<23573> A_IWL<23572> A_IWL<23571> A_IWL<23570> A_IWL<23569> A_IWL<23568> A_IWL<23567> A_IWL<23566> A_IWL<23565> A_IWL<23564> A_IWL<23563> A_IWL<23562> A_IWL<23561> A_IWL<23560> A_IWL<23559> A_IWL<23558> A_IWL<23557> A_IWL<23556> A_IWL<23555> A_IWL<23554> A_IWL<23553> A_IWL<23552> A_IWL<24575> A_IWL<24574> A_IWL<24573> A_IWL<24572> A_IWL<24571> A_IWL<24570> A_IWL<24569> A_IWL<24568> A_IWL<24567> A_IWL<24566> A_IWL<24565> A_IWL<24564> A_IWL<24563> A_IWL<24562> A_IWL<24561> A_IWL<24560> A_IWL<24559> A_IWL<24558> A_IWL<24557> A_IWL<24556> A_IWL<24555> A_IWL<24554> A_IWL<24553> A_IWL<24552> A_IWL<24551> A_IWL<24550> A_IWL<24549> A_IWL<24548> A_IWL<24547> A_IWL<24546> A_IWL<24545> A_IWL<24544> A_IWL<24543> A_IWL<24542> A_IWL<24541> A_IWL<24540> A_IWL<24539> A_IWL<24538> A_IWL<24537> A_IWL<24536> A_IWL<24535> A_IWL<24534> A_IWL<24533> A_IWL<24532> A_IWL<24531> A_IWL<24530> A_IWL<24529> A_IWL<24528> A_IWL<24527> A_IWL<24526> A_IWL<24525> A_IWL<24524> A_IWL<24523> A_IWL<24522> A_IWL<24521> A_IWL<24520> A_IWL<24519> A_IWL<24518> A_IWL<24517> A_IWL<24516> A_IWL<24515> A_IWL<24514> A_IWL<24513> A_IWL<24512> A_IWL<24511> A_IWL<24510> A_IWL<24509> A_IWL<24508> A_IWL<24507> A_IWL<24506> A_IWL<24505> A_IWL<24504> A_IWL<24503> A_IWL<24502> A_IWL<24501> A_IWL<24500> A_IWL<24499> A_IWL<24498> A_IWL<24497> A_IWL<24496> A_IWL<24495> A_IWL<24494> A_IWL<24493> A_IWL<24492> A_IWL<24491> A_IWL<24490> A_IWL<24489> A_IWL<24488> A_IWL<24487> A_IWL<24486> A_IWL<24485> A_IWL<24484> A_IWL<24483> A_IWL<24482> A_IWL<24481> A_IWL<24480> A_IWL<24479> A_IWL<24478> A_IWL<24477> A_IWL<24476> A_IWL<24475> A_IWL<24474> A_IWL<24473> A_IWL<24472> A_IWL<24471> A_IWL<24470> A_IWL<24469> A_IWL<24468> A_IWL<24467> A_IWL<24466> A_IWL<24465> A_IWL<24464> A_IWL<24463> A_IWL<24462> A_IWL<24461> A_IWL<24460> A_IWL<24459> A_IWL<24458> A_IWL<24457> A_IWL<24456> A_IWL<24455> A_IWL<24454> A_IWL<24453> A_IWL<24452> A_IWL<24451> A_IWL<24450> A_IWL<24449> A_IWL<24448> A_IWL<24447> A_IWL<24446> A_IWL<24445> A_IWL<24444> A_IWL<24443> A_IWL<24442> A_IWL<24441> A_IWL<24440> A_IWL<24439> A_IWL<24438> A_IWL<24437> A_IWL<24436> A_IWL<24435> A_IWL<24434> A_IWL<24433> A_IWL<24432> A_IWL<24431> A_IWL<24430> A_IWL<24429> A_IWL<24428> A_IWL<24427> A_IWL<24426> A_IWL<24425> A_IWL<24424> A_IWL<24423> A_IWL<24422> A_IWL<24421> A_IWL<24420> A_IWL<24419> A_IWL<24418> A_IWL<24417> A_IWL<24416> A_IWL<24415> A_IWL<24414> A_IWL<24413> A_IWL<24412> A_IWL<24411> A_IWL<24410> A_IWL<24409> A_IWL<24408> A_IWL<24407> A_IWL<24406> A_IWL<24405> A_IWL<24404> A_IWL<24403> A_IWL<24402> A_IWL<24401> A_IWL<24400> A_IWL<24399> A_IWL<24398> A_IWL<24397> A_IWL<24396> A_IWL<24395> A_IWL<24394> A_IWL<24393> A_IWL<24392> A_IWL<24391> A_IWL<24390> A_IWL<24389> A_IWL<24388> A_IWL<24387> A_IWL<24386> A_IWL<24385> A_IWL<24384> A_IWL<24383> A_IWL<24382> A_IWL<24381> A_IWL<24380> A_IWL<24379> A_IWL<24378> A_IWL<24377> A_IWL<24376> A_IWL<24375> A_IWL<24374> A_IWL<24373> A_IWL<24372> A_IWL<24371> A_IWL<24370> A_IWL<24369> A_IWL<24368> A_IWL<24367> A_IWL<24366> A_IWL<24365> A_IWL<24364> A_IWL<24363> A_IWL<24362> A_IWL<24361> A_IWL<24360> A_IWL<24359> A_IWL<24358> A_IWL<24357> A_IWL<24356> A_IWL<24355> A_IWL<24354> A_IWL<24353> A_IWL<24352> A_IWL<24351> A_IWL<24350> A_IWL<24349> A_IWL<24348> A_IWL<24347> A_IWL<24346> A_IWL<24345> A_IWL<24344> A_IWL<24343> A_IWL<24342> A_IWL<24341> A_IWL<24340> A_IWL<24339> A_IWL<24338> A_IWL<24337> A_IWL<24336> A_IWL<24335> A_IWL<24334> A_IWL<24333> A_IWL<24332> A_IWL<24331> A_IWL<24330> A_IWL<24329> A_IWL<24328> A_IWL<24327> A_IWL<24326> A_IWL<24325> A_IWL<24324> A_IWL<24323> A_IWL<24322> A_IWL<24321> A_IWL<24320> A_IWL<24319> A_IWL<24318> A_IWL<24317> A_IWL<24316> A_IWL<24315> A_IWL<24314> A_IWL<24313> A_IWL<24312> A_IWL<24311> A_IWL<24310> A_IWL<24309> A_IWL<24308> A_IWL<24307> A_IWL<24306> A_IWL<24305> A_IWL<24304> A_IWL<24303> A_IWL<24302> A_IWL<24301> A_IWL<24300> A_IWL<24299> A_IWL<24298> A_IWL<24297> A_IWL<24296> A_IWL<24295> A_IWL<24294> A_IWL<24293> A_IWL<24292> A_IWL<24291> A_IWL<24290> A_IWL<24289> A_IWL<24288> A_IWL<24287> A_IWL<24286> A_IWL<24285> A_IWL<24284> A_IWL<24283> A_IWL<24282> A_IWL<24281> A_IWL<24280> A_IWL<24279> A_IWL<24278> A_IWL<24277> A_IWL<24276> A_IWL<24275> A_IWL<24274> A_IWL<24273> A_IWL<24272> A_IWL<24271> A_IWL<24270> A_IWL<24269> A_IWL<24268> A_IWL<24267> A_IWL<24266> A_IWL<24265> A_IWL<24264> A_IWL<24263> A_IWL<24262> A_IWL<24261> A_IWL<24260> A_IWL<24259> A_IWL<24258> A_IWL<24257> A_IWL<24256> A_IWL<24255> A_IWL<24254> A_IWL<24253> A_IWL<24252> A_IWL<24251> A_IWL<24250> A_IWL<24249> A_IWL<24248> A_IWL<24247> A_IWL<24246> A_IWL<24245> A_IWL<24244> A_IWL<24243> A_IWL<24242> A_IWL<24241> A_IWL<24240> A_IWL<24239> A_IWL<24238> A_IWL<24237> A_IWL<24236> A_IWL<24235> A_IWL<24234> A_IWL<24233> A_IWL<24232> A_IWL<24231> A_IWL<24230> A_IWL<24229> A_IWL<24228> A_IWL<24227> A_IWL<24226> A_IWL<24225> A_IWL<24224> A_IWL<24223> A_IWL<24222> A_IWL<24221> A_IWL<24220> A_IWL<24219> A_IWL<24218> A_IWL<24217> A_IWL<24216> A_IWL<24215> A_IWL<24214> A_IWL<24213> A_IWL<24212> A_IWL<24211> A_IWL<24210> A_IWL<24209> A_IWL<24208> A_IWL<24207> A_IWL<24206> A_IWL<24205> A_IWL<24204> A_IWL<24203> A_IWL<24202> A_IWL<24201> A_IWL<24200> A_IWL<24199> A_IWL<24198> A_IWL<24197> A_IWL<24196> A_IWL<24195> A_IWL<24194> A_IWL<24193> A_IWL<24192> A_IWL<24191> A_IWL<24190> A_IWL<24189> A_IWL<24188> A_IWL<24187> A_IWL<24186> A_IWL<24185> A_IWL<24184> A_IWL<24183> A_IWL<24182> A_IWL<24181> A_IWL<24180> A_IWL<24179> A_IWL<24178> A_IWL<24177> A_IWL<24176> A_IWL<24175> A_IWL<24174> A_IWL<24173> A_IWL<24172> A_IWL<24171> A_IWL<24170> A_IWL<24169> A_IWL<24168> A_IWL<24167> A_IWL<24166> A_IWL<24165> A_IWL<24164> A_IWL<24163> A_IWL<24162> A_IWL<24161> A_IWL<24160> A_IWL<24159> A_IWL<24158> A_IWL<24157> A_IWL<24156> A_IWL<24155> A_IWL<24154> A_IWL<24153> A_IWL<24152> A_IWL<24151> A_IWL<24150> A_IWL<24149> A_IWL<24148> A_IWL<24147> A_IWL<24146> A_IWL<24145> A_IWL<24144> A_IWL<24143> A_IWL<24142> A_IWL<24141> A_IWL<24140> A_IWL<24139> A_IWL<24138> A_IWL<24137> A_IWL<24136> A_IWL<24135> A_IWL<24134> A_IWL<24133> A_IWL<24132> A_IWL<24131> A_IWL<24130> A_IWL<24129> A_IWL<24128> A_IWL<24127> A_IWL<24126> A_IWL<24125> A_IWL<24124> A_IWL<24123> A_IWL<24122> A_IWL<24121> A_IWL<24120> A_IWL<24119> A_IWL<24118> A_IWL<24117> A_IWL<24116> A_IWL<24115> A_IWL<24114> A_IWL<24113> A_IWL<24112> A_IWL<24111> A_IWL<24110> A_IWL<24109> A_IWL<24108> A_IWL<24107> A_IWL<24106> A_IWL<24105> A_IWL<24104> A_IWL<24103> A_IWL<24102> A_IWL<24101> A_IWL<24100> A_IWL<24099> A_IWL<24098> A_IWL<24097> A_IWL<24096> A_IWL<24095> A_IWL<24094> A_IWL<24093> A_IWL<24092> A_IWL<24091> A_IWL<24090> A_IWL<24089> A_IWL<24088> A_IWL<24087> A_IWL<24086> A_IWL<24085> A_IWL<24084> A_IWL<24083> A_IWL<24082> A_IWL<24081> A_IWL<24080> A_IWL<24079> A_IWL<24078> A_IWL<24077> A_IWL<24076> A_IWL<24075> A_IWL<24074> A_IWL<24073> A_IWL<24072> A_IWL<24071> A_IWL<24070> A_IWL<24069> A_IWL<24068> A_IWL<24067> A_IWL<24066> A_IWL<24065> A_IWL<24064> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<46> A_BLC<93> A_BLC<92> A_BLC_TOP<93> A_BLC_TOP<92> A_BLT<93> A_BLT<92> A_BLT_TOP<93> A_BLT_TOP<92> A_IWL<23551> A_IWL<23550> A_IWL<23549> A_IWL<23548> A_IWL<23547> A_IWL<23546> A_IWL<23545> A_IWL<23544> A_IWL<23543> A_IWL<23542> A_IWL<23541> A_IWL<23540> A_IWL<23539> A_IWL<23538> A_IWL<23537> A_IWL<23536> A_IWL<23535> A_IWL<23534> A_IWL<23533> A_IWL<23532> A_IWL<23531> A_IWL<23530> A_IWL<23529> A_IWL<23528> A_IWL<23527> A_IWL<23526> A_IWL<23525> A_IWL<23524> A_IWL<23523> A_IWL<23522> A_IWL<23521> A_IWL<23520> A_IWL<23519> A_IWL<23518> A_IWL<23517> A_IWL<23516> A_IWL<23515> A_IWL<23514> A_IWL<23513> A_IWL<23512> A_IWL<23511> A_IWL<23510> A_IWL<23509> A_IWL<23508> A_IWL<23507> A_IWL<23506> A_IWL<23505> A_IWL<23504> A_IWL<23503> A_IWL<23502> A_IWL<23501> A_IWL<23500> A_IWL<23499> A_IWL<23498> A_IWL<23497> A_IWL<23496> A_IWL<23495> A_IWL<23494> A_IWL<23493> A_IWL<23492> A_IWL<23491> A_IWL<23490> A_IWL<23489> A_IWL<23488> A_IWL<23487> A_IWL<23486> A_IWL<23485> A_IWL<23484> A_IWL<23483> A_IWL<23482> A_IWL<23481> A_IWL<23480> A_IWL<23479> A_IWL<23478> A_IWL<23477> A_IWL<23476> A_IWL<23475> A_IWL<23474> A_IWL<23473> A_IWL<23472> A_IWL<23471> A_IWL<23470> A_IWL<23469> A_IWL<23468> A_IWL<23467> A_IWL<23466> A_IWL<23465> A_IWL<23464> A_IWL<23463> A_IWL<23462> A_IWL<23461> A_IWL<23460> A_IWL<23459> A_IWL<23458> A_IWL<23457> A_IWL<23456> A_IWL<23455> A_IWL<23454> A_IWL<23453> A_IWL<23452> A_IWL<23451> A_IWL<23450> A_IWL<23449> A_IWL<23448> A_IWL<23447> A_IWL<23446> A_IWL<23445> A_IWL<23444> A_IWL<23443> A_IWL<23442> A_IWL<23441> A_IWL<23440> A_IWL<23439> A_IWL<23438> A_IWL<23437> A_IWL<23436> A_IWL<23435> A_IWL<23434> A_IWL<23433> A_IWL<23432> A_IWL<23431> A_IWL<23430> A_IWL<23429> A_IWL<23428> A_IWL<23427> A_IWL<23426> A_IWL<23425> A_IWL<23424> A_IWL<23423> A_IWL<23422> A_IWL<23421> A_IWL<23420> A_IWL<23419> A_IWL<23418> A_IWL<23417> A_IWL<23416> A_IWL<23415> A_IWL<23414> A_IWL<23413> A_IWL<23412> A_IWL<23411> A_IWL<23410> A_IWL<23409> A_IWL<23408> A_IWL<23407> A_IWL<23406> A_IWL<23405> A_IWL<23404> A_IWL<23403> A_IWL<23402> A_IWL<23401> A_IWL<23400> A_IWL<23399> A_IWL<23398> A_IWL<23397> A_IWL<23396> A_IWL<23395> A_IWL<23394> A_IWL<23393> A_IWL<23392> A_IWL<23391> A_IWL<23390> A_IWL<23389> A_IWL<23388> A_IWL<23387> A_IWL<23386> A_IWL<23385> A_IWL<23384> A_IWL<23383> A_IWL<23382> A_IWL<23381> A_IWL<23380> A_IWL<23379> A_IWL<23378> A_IWL<23377> A_IWL<23376> A_IWL<23375> A_IWL<23374> A_IWL<23373> A_IWL<23372> A_IWL<23371> A_IWL<23370> A_IWL<23369> A_IWL<23368> A_IWL<23367> A_IWL<23366> A_IWL<23365> A_IWL<23364> A_IWL<23363> A_IWL<23362> A_IWL<23361> A_IWL<23360> A_IWL<23359> A_IWL<23358> A_IWL<23357> A_IWL<23356> A_IWL<23355> A_IWL<23354> A_IWL<23353> A_IWL<23352> A_IWL<23351> A_IWL<23350> A_IWL<23349> A_IWL<23348> A_IWL<23347> A_IWL<23346> A_IWL<23345> A_IWL<23344> A_IWL<23343> A_IWL<23342> A_IWL<23341> A_IWL<23340> A_IWL<23339> A_IWL<23338> A_IWL<23337> A_IWL<23336> A_IWL<23335> A_IWL<23334> A_IWL<23333> A_IWL<23332> A_IWL<23331> A_IWL<23330> A_IWL<23329> A_IWL<23328> A_IWL<23327> A_IWL<23326> A_IWL<23325> A_IWL<23324> A_IWL<23323> A_IWL<23322> A_IWL<23321> A_IWL<23320> A_IWL<23319> A_IWL<23318> A_IWL<23317> A_IWL<23316> A_IWL<23315> A_IWL<23314> A_IWL<23313> A_IWL<23312> A_IWL<23311> A_IWL<23310> A_IWL<23309> A_IWL<23308> A_IWL<23307> A_IWL<23306> A_IWL<23305> A_IWL<23304> A_IWL<23303> A_IWL<23302> A_IWL<23301> A_IWL<23300> A_IWL<23299> A_IWL<23298> A_IWL<23297> A_IWL<23296> A_IWL<23295> A_IWL<23294> A_IWL<23293> A_IWL<23292> A_IWL<23291> A_IWL<23290> A_IWL<23289> A_IWL<23288> A_IWL<23287> A_IWL<23286> A_IWL<23285> A_IWL<23284> A_IWL<23283> A_IWL<23282> A_IWL<23281> A_IWL<23280> A_IWL<23279> A_IWL<23278> A_IWL<23277> A_IWL<23276> A_IWL<23275> A_IWL<23274> A_IWL<23273> A_IWL<23272> A_IWL<23271> A_IWL<23270> A_IWL<23269> A_IWL<23268> A_IWL<23267> A_IWL<23266> A_IWL<23265> A_IWL<23264> A_IWL<23263> A_IWL<23262> A_IWL<23261> A_IWL<23260> A_IWL<23259> A_IWL<23258> A_IWL<23257> A_IWL<23256> A_IWL<23255> A_IWL<23254> A_IWL<23253> A_IWL<23252> A_IWL<23251> A_IWL<23250> A_IWL<23249> A_IWL<23248> A_IWL<23247> A_IWL<23246> A_IWL<23245> A_IWL<23244> A_IWL<23243> A_IWL<23242> A_IWL<23241> A_IWL<23240> A_IWL<23239> A_IWL<23238> A_IWL<23237> A_IWL<23236> A_IWL<23235> A_IWL<23234> A_IWL<23233> A_IWL<23232> A_IWL<23231> A_IWL<23230> A_IWL<23229> A_IWL<23228> A_IWL<23227> A_IWL<23226> A_IWL<23225> A_IWL<23224> A_IWL<23223> A_IWL<23222> A_IWL<23221> A_IWL<23220> A_IWL<23219> A_IWL<23218> A_IWL<23217> A_IWL<23216> A_IWL<23215> A_IWL<23214> A_IWL<23213> A_IWL<23212> A_IWL<23211> A_IWL<23210> A_IWL<23209> A_IWL<23208> A_IWL<23207> A_IWL<23206> A_IWL<23205> A_IWL<23204> A_IWL<23203> A_IWL<23202> A_IWL<23201> A_IWL<23200> A_IWL<23199> A_IWL<23198> A_IWL<23197> A_IWL<23196> A_IWL<23195> A_IWL<23194> A_IWL<23193> A_IWL<23192> A_IWL<23191> A_IWL<23190> A_IWL<23189> A_IWL<23188> A_IWL<23187> A_IWL<23186> A_IWL<23185> A_IWL<23184> A_IWL<23183> A_IWL<23182> A_IWL<23181> A_IWL<23180> A_IWL<23179> A_IWL<23178> A_IWL<23177> A_IWL<23176> A_IWL<23175> A_IWL<23174> A_IWL<23173> A_IWL<23172> A_IWL<23171> A_IWL<23170> A_IWL<23169> A_IWL<23168> A_IWL<23167> A_IWL<23166> A_IWL<23165> A_IWL<23164> A_IWL<23163> A_IWL<23162> A_IWL<23161> A_IWL<23160> A_IWL<23159> A_IWL<23158> A_IWL<23157> A_IWL<23156> A_IWL<23155> A_IWL<23154> A_IWL<23153> A_IWL<23152> A_IWL<23151> A_IWL<23150> A_IWL<23149> A_IWL<23148> A_IWL<23147> A_IWL<23146> A_IWL<23145> A_IWL<23144> A_IWL<23143> A_IWL<23142> A_IWL<23141> A_IWL<23140> A_IWL<23139> A_IWL<23138> A_IWL<23137> A_IWL<23136> A_IWL<23135> A_IWL<23134> A_IWL<23133> A_IWL<23132> A_IWL<23131> A_IWL<23130> A_IWL<23129> A_IWL<23128> A_IWL<23127> A_IWL<23126> A_IWL<23125> A_IWL<23124> A_IWL<23123> A_IWL<23122> A_IWL<23121> A_IWL<23120> A_IWL<23119> A_IWL<23118> A_IWL<23117> A_IWL<23116> A_IWL<23115> A_IWL<23114> A_IWL<23113> A_IWL<23112> A_IWL<23111> A_IWL<23110> A_IWL<23109> A_IWL<23108> A_IWL<23107> A_IWL<23106> A_IWL<23105> A_IWL<23104> A_IWL<23103> A_IWL<23102> A_IWL<23101> A_IWL<23100> A_IWL<23099> A_IWL<23098> A_IWL<23097> A_IWL<23096> A_IWL<23095> A_IWL<23094> A_IWL<23093> A_IWL<23092> A_IWL<23091> A_IWL<23090> A_IWL<23089> A_IWL<23088> A_IWL<23087> A_IWL<23086> A_IWL<23085> A_IWL<23084> A_IWL<23083> A_IWL<23082> A_IWL<23081> A_IWL<23080> A_IWL<23079> A_IWL<23078> A_IWL<23077> A_IWL<23076> A_IWL<23075> A_IWL<23074> A_IWL<23073> A_IWL<23072> A_IWL<23071> A_IWL<23070> A_IWL<23069> A_IWL<23068> A_IWL<23067> A_IWL<23066> A_IWL<23065> A_IWL<23064> A_IWL<23063> A_IWL<23062> A_IWL<23061> A_IWL<23060> A_IWL<23059> A_IWL<23058> A_IWL<23057> A_IWL<23056> A_IWL<23055> A_IWL<23054> A_IWL<23053> A_IWL<23052> A_IWL<23051> A_IWL<23050> A_IWL<23049> A_IWL<23048> A_IWL<23047> A_IWL<23046> A_IWL<23045> A_IWL<23044> A_IWL<23043> A_IWL<23042> A_IWL<23041> A_IWL<23040> A_IWL<24063> A_IWL<24062> A_IWL<24061> A_IWL<24060> A_IWL<24059> A_IWL<24058> A_IWL<24057> A_IWL<24056> A_IWL<24055> A_IWL<24054> A_IWL<24053> A_IWL<24052> A_IWL<24051> A_IWL<24050> A_IWL<24049> A_IWL<24048> A_IWL<24047> A_IWL<24046> A_IWL<24045> A_IWL<24044> A_IWL<24043> A_IWL<24042> A_IWL<24041> A_IWL<24040> A_IWL<24039> A_IWL<24038> A_IWL<24037> A_IWL<24036> A_IWL<24035> A_IWL<24034> A_IWL<24033> A_IWL<24032> A_IWL<24031> A_IWL<24030> A_IWL<24029> A_IWL<24028> A_IWL<24027> A_IWL<24026> A_IWL<24025> A_IWL<24024> A_IWL<24023> A_IWL<24022> A_IWL<24021> A_IWL<24020> A_IWL<24019> A_IWL<24018> A_IWL<24017> A_IWL<24016> A_IWL<24015> A_IWL<24014> A_IWL<24013> A_IWL<24012> A_IWL<24011> A_IWL<24010> A_IWL<24009> A_IWL<24008> A_IWL<24007> A_IWL<24006> A_IWL<24005> A_IWL<24004> A_IWL<24003> A_IWL<24002> A_IWL<24001> A_IWL<24000> A_IWL<23999> A_IWL<23998> A_IWL<23997> A_IWL<23996> A_IWL<23995> A_IWL<23994> A_IWL<23993> A_IWL<23992> A_IWL<23991> A_IWL<23990> A_IWL<23989> A_IWL<23988> A_IWL<23987> A_IWL<23986> A_IWL<23985> A_IWL<23984> A_IWL<23983> A_IWL<23982> A_IWL<23981> A_IWL<23980> A_IWL<23979> A_IWL<23978> A_IWL<23977> A_IWL<23976> A_IWL<23975> A_IWL<23974> A_IWL<23973> A_IWL<23972> A_IWL<23971> A_IWL<23970> A_IWL<23969> A_IWL<23968> A_IWL<23967> A_IWL<23966> A_IWL<23965> A_IWL<23964> A_IWL<23963> A_IWL<23962> A_IWL<23961> A_IWL<23960> A_IWL<23959> A_IWL<23958> A_IWL<23957> A_IWL<23956> A_IWL<23955> A_IWL<23954> A_IWL<23953> A_IWL<23952> A_IWL<23951> A_IWL<23950> A_IWL<23949> A_IWL<23948> A_IWL<23947> A_IWL<23946> A_IWL<23945> A_IWL<23944> A_IWL<23943> A_IWL<23942> A_IWL<23941> A_IWL<23940> A_IWL<23939> A_IWL<23938> A_IWL<23937> A_IWL<23936> A_IWL<23935> A_IWL<23934> A_IWL<23933> A_IWL<23932> A_IWL<23931> A_IWL<23930> A_IWL<23929> A_IWL<23928> A_IWL<23927> A_IWL<23926> A_IWL<23925> A_IWL<23924> A_IWL<23923> A_IWL<23922> A_IWL<23921> A_IWL<23920> A_IWL<23919> A_IWL<23918> A_IWL<23917> A_IWL<23916> A_IWL<23915> A_IWL<23914> A_IWL<23913> A_IWL<23912> A_IWL<23911> A_IWL<23910> A_IWL<23909> A_IWL<23908> A_IWL<23907> A_IWL<23906> A_IWL<23905> A_IWL<23904> A_IWL<23903> A_IWL<23902> A_IWL<23901> A_IWL<23900> A_IWL<23899> A_IWL<23898> A_IWL<23897> A_IWL<23896> A_IWL<23895> A_IWL<23894> A_IWL<23893> A_IWL<23892> A_IWL<23891> A_IWL<23890> A_IWL<23889> A_IWL<23888> A_IWL<23887> A_IWL<23886> A_IWL<23885> A_IWL<23884> A_IWL<23883> A_IWL<23882> A_IWL<23881> A_IWL<23880> A_IWL<23879> A_IWL<23878> A_IWL<23877> A_IWL<23876> A_IWL<23875> A_IWL<23874> A_IWL<23873> A_IWL<23872> A_IWL<23871> A_IWL<23870> A_IWL<23869> A_IWL<23868> A_IWL<23867> A_IWL<23866> A_IWL<23865> A_IWL<23864> A_IWL<23863> A_IWL<23862> A_IWL<23861> A_IWL<23860> A_IWL<23859> A_IWL<23858> A_IWL<23857> A_IWL<23856> A_IWL<23855> A_IWL<23854> A_IWL<23853> A_IWL<23852> A_IWL<23851> A_IWL<23850> A_IWL<23849> A_IWL<23848> A_IWL<23847> A_IWL<23846> A_IWL<23845> A_IWL<23844> A_IWL<23843> A_IWL<23842> A_IWL<23841> A_IWL<23840> A_IWL<23839> A_IWL<23838> A_IWL<23837> A_IWL<23836> A_IWL<23835> A_IWL<23834> A_IWL<23833> A_IWL<23832> A_IWL<23831> A_IWL<23830> A_IWL<23829> A_IWL<23828> A_IWL<23827> A_IWL<23826> A_IWL<23825> A_IWL<23824> A_IWL<23823> A_IWL<23822> A_IWL<23821> A_IWL<23820> A_IWL<23819> A_IWL<23818> A_IWL<23817> A_IWL<23816> A_IWL<23815> A_IWL<23814> A_IWL<23813> A_IWL<23812> A_IWL<23811> A_IWL<23810> A_IWL<23809> A_IWL<23808> A_IWL<23807> A_IWL<23806> A_IWL<23805> A_IWL<23804> A_IWL<23803> A_IWL<23802> A_IWL<23801> A_IWL<23800> A_IWL<23799> A_IWL<23798> A_IWL<23797> A_IWL<23796> A_IWL<23795> A_IWL<23794> A_IWL<23793> A_IWL<23792> A_IWL<23791> A_IWL<23790> A_IWL<23789> A_IWL<23788> A_IWL<23787> A_IWL<23786> A_IWL<23785> A_IWL<23784> A_IWL<23783> A_IWL<23782> A_IWL<23781> A_IWL<23780> A_IWL<23779> A_IWL<23778> A_IWL<23777> A_IWL<23776> A_IWL<23775> A_IWL<23774> A_IWL<23773> A_IWL<23772> A_IWL<23771> A_IWL<23770> A_IWL<23769> A_IWL<23768> A_IWL<23767> A_IWL<23766> A_IWL<23765> A_IWL<23764> A_IWL<23763> A_IWL<23762> A_IWL<23761> A_IWL<23760> A_IWL<23759> A_IWL<23758> A_IWL<23757> A_IWL<23756> A_IWL<23755> A_IWL<23754> A_IWL<23753> A_IWL<23752> A_IWL<23751> A_IWL<23750> A_IWL<23749> A_IWL<23748> A_IWL<23747> A_IWL<23746> A_IWL<23745> A_IWL<23744> A_IWL<23743> A_IWL<23742> A_IWL<23741> A_IWL<23740> A_IWL<23739> A_IWL<23738> A_IWL<23737> A_IWL<23736> A_IWL<23735> A_IWL<23734> A_IWL<23733> A_IWL<23732> A_IWL<23731> A_IWL<23730> A_IWL<23729> A_IWL<23728> A_IWL<23727> A_IWL<23726> A_IWL<23725> A_IWL<23724> A_IWL<23723> A_IWL<23722> A_IWL<23721> A_IWL<23720> A_IWL<23719> A_IWL<23718> A_IWL<23717> A_IWL<23716> A_IWL<23715> A_IWL<23714> A_IWL<23713> A_IWL<23712> A_IWL<23711> A_IWL<23710> A_IWL<23709> A_IWL<23708> A_IWL<23707> A_IWL<23706> A_IWL<23705> A_IWL<23704> A_IWL<23703> A_IWL<23702> A_IWL<23701> A_IWL<23700> A_IWL<23699> A_IWL<23698> A_IWL<23697> A_IWL<23696> A_IWL<23695> A_IWL<23694> A_IWL<23693> A_IWL<23692> A_IWL<23691> A_IWL<23690> A_IWL<23689> A_IWL<23688> A_IWL<23687> A_IWL<23686> A_IWL<23685> A_IWL<23684> A_IWL<23683> A_IWL<23682> A_IWL<23681> A_IWL<23680> A_IWL<23679> A_IWL<23678> A_IWL<23677> A_IWL<23676> A_IWL<23675> A_IWL<23674> A_IWL<23673> A_IWL<23672> A_IWL<23671> A_IWL<23670> A_IWL<23669> A_IWL<23668> A_IWL<23667> A_IWL<23666> A_IWL<23665> A_IWL<23664> A_IWL<23663> A_IWL<23662> A_IWL<23661> A_IWL<23660> A_IWL<23659> A_IWL<23658> A_IWL<23657> A_IWL<23656> A_IWL<23655> A_IWL<23654> A_IWL<23653> A_IWL<23652> A_IWL<23651> A_IWL<23650> A_IWL<23649> A_IWL<23648> A_IWL<23647> A_IWL<23646> A_IWL<23645> A_IWL<23644> A_IWL<23643> A_IWL<23642> A_IWL<23641> A_IWL<23640> A_IWL<23639> A_IWL<23638> A_IWL<23637> A_IWL<23636> A_IWL<23635> A_IWL<23634> A_IWL<23633> A_IWL<23632> A_IWL<23631> A_IWL<23630> A_IWL<23629> A_IWL<23628> A_IWL<23627> A_IWL<23626> A_IWL<23625> A_IWL<23624> A_IWL<23623> A_IWL<23622> A_IWL<23621> A_IWL<23620> A_IWL<23619> A_IWL<23618> A_IWL<23617> A_IWL<23616> A_IWL<23615> A_IWL<23614> A_IWL<23613> A_IWL<23612> A_IWL<23611> A_IWL<23610> A_IWL<23609> A_IWL<23608> A_IWL<23607> A_IWL<23606> A_IWL<23605> A_IWL<23604> A_IWL<23603> A_IWL<23602> A_IWL<23601> A_IWL<23600> A_IWL<23599> A_IWL<23598> A_IWL<23597> A_IWL<23596> A_IWL<23595> A_IWL<23594> A_IWL<23593> A_IWL<23592> A_IWL<23591> A_IWL<23590> A_IWL<23589> A_IWL<23588> A_IWL<23587> A_IWL<23586> A_IWL<23585> A_IWL<23584> A_IWL<23583> A_IWL<23582> A_IWL<23581> A_IWL<23580> A_IWL<23579> A_IWL<23578> A_IWL<23577> A_IWL<23576> A_IWL<23575> A_IWL<23574> A_IWL<23573> A_IWL<23572> A_IWL<23571> A_IWL<23570> A_IWL<23569> A_IWL<23568> A_IWL<23567> A_IWL<23566> A_IWL<23565> A_IWL<23564> A_IWL<23563> A_IWL<23562> A_IWL<23561> A_IWL<23560> A_IWL<23559> A_IWL<23558> A_IWL<23557> A_IWL<23556> A_IWL<23555> A_IWL<23554> A_IWL<23553> A_IWL<23552> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<45> A_BLC<91> A_BLC<90> A_BLC_TOP<91> A_BLC_TOP<90> A_BLT<91> A_BLT<90> A_BLT_TOP<91> A_BLT_TOP<90> A_IWL<23039> A_IWL<23038> A_IWL<23037> A_IWL<23036> A_IWL<23035> A_IWL<23034> A_IWL<23033> A_IWL<23032> A_IWL<23031> A_IWL<23030> A_IWL<23029> A_IWL<23028> A_IWL<23027> A_IWL<23026> A_IWL<23025> A_IWL<23024> A_IWL<23023> A_IWL<23022> A_IWL<23021> A_IWL<23020> A_IWL<23019> A_IWL<23018> A_IWL<23017> A_IWL<23016> A_IWL<23015> A_IWL<23014> A_IWL<23013> A_IWL<23012> A_IWL<23011> A_IWL<23010> A_IWL<23009> A_IWL<23008> A_IWL<23007> A_IWL<23006> A_IWL<23005> A_IWL<23004> A_IWL<23003> A_IWL<23002> A_IWL<23001> A_IWL<23000> A_IWL<22999> A_IWL<22998> A_IWL<22997> A_IWL<22996> A_IWL<22995> A_IWL<22994> A_IWL<22993> A_IWL<22992> A_IWL<22991> A_IWL<22990> A_IWL<22989> A_IWL<22988> A_IWL<22987> A_IWL<22986> A_IWL<22985> A_IWL<22984> A_IWL<22983> A_IWL<22982> A_IWL<22981> A_IWL<22980> A_IWL<22979> A_IWL<22978> A_IWL<22977> A_IWL<22976> A_IWL<22975> A_IWL<22974> A_IWL<22973> A_IWL<22972> A_IWL<22971> A_IWL<22970> A_IWL<22969> A_IWL<22968> A_IWL<22967> A_IWL<22966> A_IWL<22965> A_IWL<22964> A_IWL<22963> A_IWL<22962> A_IWL<22961> A_IWL<22960> A_IWL<22959> A_IWL<22958> A_IWL<22957> A_IWL<22956> A_IWL<22955> A_IWL<22954> A_IWL<22953> A_IWL<22952> A_IWL<22951> A_IWL<22950> A_IWL<22949> A_IWL<22948> A_IWL<22947> A_IWL<22946> A_IWL<22945> A_IWL<22944> A_IWL<22943> A_IWL<22942> A_IWL<22941> A_IWL<22940> A_IWL<22939> A_IWL<22938> A_IWL<22937> A_IWL<22936> A_IWL<22935> A_IWL<22934> A_IWL<22933> A_IWL<22932> A_IWL<22931> A_IWL<22930> A_IWL<22929> A_IWL<22928> A_IWL<22927> A_IWL<22926> A_IWL<22925> A_IWL<22924> A_IWL<22923> A_IWL<22922> A_IWL<22921> A_IWL<22920> A_IWL<22919> A_IWL<22918> A_IWL<22917> A_IWL<22916> A_IWL<22915> A_IWL<22914> A_IWL<22913> A_IWL<22912> A_IWL<22911> A_IWL<22910> A_IWL<22909> A_IWL<22908> A_IWL<22907> A_IWL<22906> A_IWL<22905> A_IWL<22904> A_IWL<22903> A_IWL<22902> A_IWL<22901> A_IWL<22900> A_IWL<22899> A_IWL<22898> A_IWL<22897> A_IWL<22896> A_IWL<22895> A_IWL<22894> A_IWL<22893> A_IWL<22892> A_IWL<22891> A_IWL<22890> A_IWL<22889> A_IWL<22888> A_IWL<22887> A_IWL<22886> A_IWL<22885> A_IWL<22884> A_IWL<22883> A_IWL<22882> A_IWL<22881> A_IWL<22880> A_IWL<22879> A_IWL<22878> A_IWL<22877> A_IWL<22876> A_IWL<22875> A_IWL<22874> A_IWL<22873> A_IWL<22872> A_IWL<22871> A_IWL<22870> A_IWL<22869> A_IWL<22868> A_IWL<22867> A_IWL<22866> A_IWL<22865> A_IWL<22864> A_IWL<22863> A_IWL<22862> A_IWL<22861> A_IWL<22860> A_IWL<22859> A_IWL<22858> A_IWL<22857> A_IWL<22856> A_IWL<22855> A_IWL<22854> A_IWL<22853> A_IWL<22852> A_IWL<22851> A_IWL<22850> A_IWL<22849> A_IWL<22848> A_IWL<22847> A_IWL<22846> A_IWL<22845> A_IWL<22844> A_IWL<22843> A_IWL<22842> A_IWL<22841> A_IWL<22840> A_IWL<22839> A_IWL<22838> A_IWL<22837> A_IWL<22836> A_IWL<22835> A_IWL<22834> A_IWL<22833> A_IWL<22832> A_IWL<22831> A_IWL<22830> A_IWL<22829> A_IWL<22828> A_IWL<22827> A_IWL<22826> A_IWL<22825> A_IWL<22824> A_IWL<22823> A_IWL<22822> A_IWL<22821> A_IWL<22820> A_IWL<22819> A_IWL<22818> A_IWL<22817> A_IWL<22816> A_IWL<22815> A_IWL<22814> A_IWL<22813> A_IWL<22812> A_IWL<22811> A_IWL<22810> A_IWL<22809> A_IWL<22808> A_IWL<22807> A_IWL<22806> A_IWL<22805> A_IWL<22804> A_IWL<22803> A_IWL<22802> A_IWL<22801> A_IWL<22800> A_IWL<22799> A_IWL<22798> A_IWL<22797> A_IWL<22796> A_IWL<22795> A_IWL<22794> A_IWL<22793> A_IWL<22792> A_IWL<22791> A_IWL<22790> A_IWL<22789> A_IWL<22788> A_IWL<22787> A_IWL<22786> A_IWL<22785> A_IWL<22784> A_IWL<22783> A_IWL<22782> A_IWL<22781> A_IWL<22780> A_IWL<22779> A_IWL<22778> A_IWL<22777> A_IWL<22776> A_IWL<22775> A_IWL<22774> A_IWL<22773> A_IWL<22772> A_IWL<22771> A_IWL<22770> A_IWL<22769> A_IWL<22768> A_IWL<22767> A_IWL<22766> A_IWL<22765> A_IWL<22764> A_IWL<22763> A_IWL<22762> A_IWL<22761> A_IWL<22760> A_IWL<22759> A_IWL<22758> A_IWL<22757> A_IWL<22756> A_IWL<22755> A_IWL<22754> A_IWL<22753> A_IWL<22752> A_IWL<22751> A_IWL<22750> A_IWL<22749> A_IWL<22748> A_IWL<22747> A_IWL<22746> A_IWL<22745> A_IWL<22744> A_IWL<22743> A_IWL<22742> A_IWL<22741> A_IWL<22740> A_IWL<22739> A_IWL<22738> A_IWL<22737> A_IWL<22736> A_IWL<22735> A_IWL<22734> A_IWL<22733> A_IWL<22732> A_IWL<22731> A_IWL<22730> A_IWL<22729> A_IWL<22728> A_IWL<22727> A_IWL<22726> A_IWL<22725> A_IWL<22724> A_IWL<22723> A_IWL<22722> A_IWL<22721> A_IWL<22720> A_IWL<22719> A_IWL<22718> A_IWL<22717> A_IWL<22716> A_IWL<22715> A_IWL<22714> A_IWL<22713> A_IWL<22712> A_IWL<22711> A_IWL<22710> A_IWL<22709> A_IWL<22708> A_IWL<22707> A_IWL<22706> A_IWL<22705> A_IWL<22704> A_IWL<22703> A_IWL<22702> A_IWL<22701> A_IWL<22700> A_IWL<22699> A_IWL<22698> A_IWL<22697> A_IWL<22696> A_IWL<22695> A_IWL<22694> A_IWL<22693> A_IWL<22692> A_IWL<22691> A_IWL<22690> A_IWL<22689> A_IWL<22688> A_IWL<22687> A_IWL<22686> A_IWL<22685> A_IWL<22684> A_IWL<22683> A_IWL<22682> A_IWL<22681> A_IWL<22680> A_IWL<22679> A_IWL<22678> A_IWL<22677> A_IWL<22676> A_IWL<22675> A_IWL<22674> A_IWL<22673> A_IWL<22672> A_IWL<22671> A_IWL<22670> A_IWL<22669> A_IWL<22668> A_IWL<22667> A_IWL<22666> A_IWL<22665> A_IWL<22664> A_IWL<22663> A_IWL<22662> A_IWL<22661> A_IWL<22660> A_IWL<22659> A_IWL<22658> A_IWL<22657> A_IWL<22656> A_IWL<22655> A_IWL<22654> A_IWL<22653> A_IWL<22652> A_IWL<22651> A_IWL<22650> A_IWL<22649> A_IWL<22648> A_IWL<22647> A_IWL<22646> A_IWL<22645> A_IWL<22644> A_IWL<22643> A_IWL<22642> A_IWL<22641> A_IWL<22640> A_IWL<22639> A_IWL<22638> A_IWL<22637> A_IWL<22636> A_IWL<22635> A_IWL<22634> A_IWL<22633> A_IWL<22632> A_IWL<22631> A_IWL<22630> A_IWL<22629> A_IWL<22628> A_IWL<22627> A_IWL<22626> A_IWL<22625> A_IWL<22624> A_IWL<22623> A_IWL<22622> A_IWL<22621> A_IWL<22620> A_IWL<22619> A_IWL<22618> A_IWL<22617> A_IWL<22616> A_IWL<22615> A_IWL<22614> A_IWL<22613> A_IWL<22612> A_IWL<22611> A_IWL<22610> A_IWL<22609> A_IWL<22608> A_IWL<22607> A_IWL<22606> A_IWL<22605> A_IWL<22604> A_IWL<22603> A_IWL<22602> A_IWL<22601> A_IWL<22600> A_IWL<22599> A_IWL<22598> A_IWL<22597> A_IWL<22596> A_IWL<22595> A_IWL<22594> A_IWL<22593> A_IWL<22592> A_IWL<22591> A_IWL<22590> A_IWL<22589> A_IWL<22588> A_IWL<22587> A_IWL<22586> A_IWL<22585> A_IWL<22584> A_IWL<22583> A_IWL<22582> A_IWL<22581> A_IWL<22580> A_IWL<22579> A_IWL<22578> A_IWL<22577> A_IWL<22576> A_IWL<22575> A_IWL<22574> A_IWL<22573> A_IWL<22572> A_IWL<22571> A_IWL<22570> A_IWL<22569> A_IWL<22568> A_IWL<22567> A_IWL<22566> A_IWL<22565> A_IWL<22564> A_IWL<22563> A_IWL<22562> A_IWL<22561> A_IWL<22560> A_IWL<22559> A_IWL<22558> A_IWL<22557> A_IWL<22556> A_IWL<22555> A_IWL<22554> A_IWL<22553> A_IWL<22552> A_IWL<22551> A_IWL<22550> A_IWL<22549> A_IWL<22548> A_IWL<22547> A_IWL<22546> A_IWL<22545> A_IWL<22544> A_IWL<22543> A_IWL<22542> A_IWL<22541> A_IWL<22540> A_IWL<22539> A_IWL<22538> A_IWL<22537> A_IWL<22536> A_IWL<22535> A_IWL<22534> A_IWL<22533> A_IWL<22532> A_IWL<22531> A_IWL<22530> A_IWL<22529> A_IWL<22528> A_IWL<23551> A_IWL<23550> A_IWL<23549> A_IWL<23548> A_IWL<23547> A_IWL<23546> A_IWL<23545> A_IWL<23544> A_IWL<23543> A_IWL<23542> A_IWL<23541> A_IWL<23540> A_IWL<23539> A_IWL<23538> A_IWL<23537> A_IWL<23536> A_IWL<23535> A_IWL<23534> A_IWL<23533> A_IWL<23532> A_IWL<23531> A_IWL<23530> A_IWL<23529> A_IWL<23528> A_IWL<23527> A_IWL<23526> A_IWL<23525> A_IWL<23524> A_IWL<23523> A_IWL<23522> A_IWL<23521> A_IWL<23520> A_IWL<23519> A_IWL<23518> A_IWL<23517> A_IWL<23516> A_IWL<23515> A_IWL<23514> A_IWL<23513> A_IWL<23512> A_IWL<23511> A_IWL<23510> A_IWL<23509> A_IWL<23508> A_IWL<23507> A_IWL<23506> A_IWL<23505> A_IWL<23504> A_IWL<23503> A_IWL<23502> A_IWL<23501> A_IWL<23500> A_IWL<23499> A_IWL<23498> A_IWL<23497> A_IWL<23496> A_IWL<23495> A_IWL<23494> A_IWL<23493> A_IWL<23492> A_IWL<23491> A_IWL<23490> A_IWL<23489> A_IWL<23488> A_IWL<23487> A_IWL<23486> A_IWL<23485> A_IWL<23484> A_IWL<23483> A_IWL<23482> A_IWL<23481> A_IWL<23480> A_IWL<23479> A_IWL<23478> A_IWL<23477> A_IWL<23476> A_IWL<23475> A_IWL<23474> A_IWL<23473> A_IWL<23472> A_IWL<23471> A_IWL<23470> A_IWL<23469> A_IWL<23468> A_IWL<23467> A_IWL<23466> A_IWL<23465> A_IWL<23464> A_IWL<23463> A_IWL<23462> A_IWL<23461> A_IWL<23460> A_IWL<23459> A_IWL<23458> A_IWL<23457> A_IWL<23456> A_IWL<23455> A_IWL<23454> A_IWL<23453> A_IWL<23452> A_IWL<23451> A_IWL<23450> A_IWL<23449> A_IWL<23448> A_IWL<23447> A_IWL<23446> A_IWL<23445> A_IWL<23444> A_IWL<23443> A_IWL<23442> A_IWL<23441> A_IWL<23440> A_IWL<23439> A_IWL<23438> A_IWL<23437> A_IWL<23436> A_IWL<23435> A_IWL<23434> A_IWL<23433> A_IWL<23432> A_IWL<23431> A_IWL<23430> A_IWL<23429> A_IWL<23428> A_IWL<23427> A_IWL<23426> A_IWL<23425> A_IWL<23424> A_IWL<23423> A_IWL<23422> A_IWL<23421> A_IWL<23420> A_IWL<23419> A_IWL<23418> A_IWL<23417> A_IWL<23416> A_IWL<23415> A_IWL<23414> A_IWL<23413> A_IWL<23412> A_IWL<23411> A_IWL<23410> A_IWL<23409> A_IWL<23408> A_IWL<23407> A_IWL<23406> A_IWL<23405> A_IWL<23404> A_IWL<23403> A_IWL<23402> A_IWL<23401> A_IWL<23400> A_IWL<23399> A_IWL<23398> A_IWL<23397> A_IWL<23396> A_IWL<23395> A_IWL<23394> A_IWL<23393> A_IWL<23392> A_IWL<23391> A_IWL<23390> A_IWL<23389> A_IWL<23388> A_IWL<23387> A_IWL<23386> A_IWL<23385> A_IWL<23384> A_IWL<23383> A_IWL<23382> A_IWL<23381> A_IWL<23380> A_IWL<23379> A_IWL<23378> A_IWL<23377> A_IWL<23376> A_IWL<23375> A_IWL<23374> A_IWL<23373> A_IWL<23372> A_IWL<23371> A_IWL<23370> A_IWL<23369> A_IWL<23368> A_IWL<23367> A_IWL<23366> A_IWL<23365> A_IWL<23364> A_IWL<23363> A_IWL<23362> A_IWL<23361> A_IWL<23360> A_IWL<23359> A_IWL<23358> A_IWL<23357> A_IWL<23356> A_IWL<23355> A_IWL<23354> A_IWL<23353> A_IWL<23352> A_IWL<23351> A_IWL<23350> A_IWL<23349> A_IWL<23348> A_IWL<23347> A_IWL<23346> A_IWL<23345> A_IWL<23344> A_IWL<23343> A_IWL<23342> A_IWL<23341> A_IWL<23340> A_IWL<23339> A_IWL<23338> A_IWL<23337> A_IWL<23336> A_IWL<23335> A_IWL<23334> A_IWL<23333> A_IWL<23332> A_IWL<23331> A_IWL<23330> A_IWL<23329> A_IWL<23328> A_IWL<23327> A_IWL<23326> A_IWL<23325> A_IWL<23324> A_IWL<23323> A_IWL<23322> A_IWL<23321> A_IWL<23320> A_IWL<23319> A_IWL<23318> A_IWL<23317> A_IWL<23316> A_IWL<23315> A_IWL<23314> A_IWL<23313> A_IWL<23312> A_IWL<23311> A_IWL<23310> A_IWL<23309> A_IWL<23308> A_IWL<23307> A_IWL<23306> A_IWL<23305> A_IWL<23304> A_IWL<23303> A_IWL<23302> A_IWL<23301> A_IWL<23300> A_IWL<23299> A_IWL<23298> A_IWL<23297> A_IWL<23296> A_IWL<23295> A_IWL<23294> A_IWL<23293> A_IWL<23292> A_IWL<23291> A_IWL<23290> A_IWL<23289> A_IWL<23288> A_IWL<23287> A_IWL<23286> A_IWL<23285> A_IWL<23284> A_IWL<23283> A_IWL<23282> A_IWL<23281> A_IWL<23280> A_IWL<23279> A_IWL<23278> A_IWL<23277> A_IWL<23276> A_IWL<23275> A_IWL<23274> A_IWL<23273> A_IWL<23272> A_IWL<23271> A_IWL<23270> A_IWL<23269> A_IWL<23268> A_IWL<23267> A_IWL<23266> A_IWL<23265> A_IWL<23264> A_IWL<23263> A_IWL<23262> A_IWL<23261> A_IWL<23260> A_IWL<23259> A_IWL<23258> A_IWL<23257> A_IWL<23256> A_IWL<23255> A_IWL<23254> A_IWL<23253> A_IWL<23252> A_IWL<23251> A_IWL<23250> A_IWL<23249> A_IWL<23248> A_IWL<23247> A_IWL<23246> A_IWL<23245> A_IWL<23244> A_IWL<23243> A_IWL<23242> A_IWL<23241> A_IWL<23240> A_IWL<23239> A_IWL<23238> A_IWL<23237> A_IWL<23236> A_IWL<23235> A_IWL<23234> A_IWL<23233> A_IWL<23232> A_IWL<23231> A_IWL<23230> A_IWL<23229> A_IWL<23228> A_IWL<23227> A_IWL<23226> A_IWL<23225> A_IWL<23224> A_IWL<23223> A_IWL<23222> A_IWL<23221> A_IWL<23220> A_IWL<23219> A_IWL<23218> A_IWL<23217> A_IWL<23216> A_IWL<23215> A_IWL<23214> A_IWL<23213> A_IWL<23212> A_IWL<23211> A_IWL<23210> A_IWL<23209> A_IWL<23208> A_IWL<23207> A_IWL<23206> A_IWL<23205> A_IWL<23204> A_IWL<23203> A_IWL<23202> A_IWL<23201> A_IWL<23200> A_IWL<23199> A_IWL<23198> A_IWL<23197> A_IWL<23196> A_IWL<23195> A_IWL<23194> A_IWL<23193> A_IWL<23192> A_IWL<23191> A_IWL<23190> A_IWL<23189> A_IWL<23188> A_IWL<23187> A_IWL<23186> A_IWL<23185> A_IWL<23184> A_IWL<23183> A_IWL<23182> A_IWL<23181> A_IWL<23180> A_IWL<23179> A_IWL<23178> A_IWL<23177> A_IWL<23176> A_IWL<23175> A_IWL<23174> A_IWL<23173> A_IWL<23172> A_IWL<23171> A_IWL<23170> A_IWL<23169> A_IWL<23168> A_IWL<23167> A_IWL<23166> A_IWL<23165> A_IWL<23164> A_IWL<23163> A_IWL<23162> A_IWL<23161> A_IWL<23160> A_IWL<23159> A_IWL<23158> A_IWL<23157> A_IWL<23156> A_IWL<23155> A_IWL<23154> A_IWL<23153> A_IWL<23152> A_IWL<23151> A_IWL<23150> A_IWL<23149> A_IWL<23148> A_IWL<23147> A_IWL<23146> A_IWL<23145> A_IWL<23144> A_IWL<23143> A_IWL<23142> A_IWL<23141> A_IWL<23140> A_IWL<23139> A_IWL<23138> A_IWL<23137> A_IWL<23136> A_IWL<23135> A_IWL<23134> A_IWL<23133> A_IWL<23132> A_IWL<23131> A_IWL<23130> A_IWL<23129> A_IWL<23128> A_IWL<23127> A_IWL<23126> A_IWL<23125> A_IWL<23124> A_IWL<23123> A_IWL<23122> A_IWL<23121> A_IWL<23120> A_IWL<23119> A_IWL<23118> A_IWL<23117> A_IWL<23116> A_IWL<23115> A_IWL<23114> A_IWL<23113> A_IWL<23112> A_IWL<23111> A_IWL<23110> A_IWL<23109> A_IWL<23108> A_IWL<23107> A_IWL<23106> A_IWL<23105> A_IWL<23104> A_IWL<23103> A_IWL<23102> A_IWL<23101> A_IWL<23100> A_IWL<23099> A_IWL<23098> A_IWL<23097> A_IWL<23096> A_IWL<23095> A_IWL<23094> A_IWL<23093> A_IWL<23092> A_IWL<23091> A_IWL<23090> A_IWL<23089> A_IWL<23088> A_IWL<23087> A_IWL<23086> A_IWL<23085> A_IWL<23084> A_IWL<23083> A_IWL<23082> A_IWL<23081> A_IWL<23080> A_IWL<23079> A_IWL<23078> A_IWL<23077> A_IWL<23076> A_IWL<23075> A_IWL<23074> A_IWL<23073> A_IWL<23072> A_IWL<23071> A_IWL<23070> A_IWL<23069> A_IWL<23068> A_IWL<23067> A_IWL<23066> A_IWL<23065> A_IWL<23064> A_IWL<23063> A_IWL<23062> A_IWL<23061> A_IWL<23060> A_IWL<23059> A_IWL<23058> A_IWL<23057> A_IWL<23056> A_IWL<23055> A_IWL<23054> A_IWL<23053> A_IWL<23052> A_IWL<23051> A_IWL<23050> A_IWL<23049> A_IWL<23048> A_IWL<23047> A_IWL<23046> A_IWL<23045> A_IWL<23044> A_IWL<23043> A_IWL<23042> A_IWL<23041> A_IWL<23040> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<44> A_BLC<89> A_BLC<88> A_BLC_TOP<89> A_BLC_TOP<88> A_BLT<89> A_BLT<88> A_BLT_TOP<89> A_BLT_TOP<88> A_IWL<22527> A_IWL<22526> A_IWL<22525> A_IWL<22524> A_IWL<22523> A_IWL<22522> A_IWL<22521> A_IWL<22520> A_IWL<22519> A_IWL<22518> A_IWL<22517> A_IWL<22516> A_IWL<22515> A_IWL<22514> A_IWL<22513> A_IWL<22512> A_IWL<22511> A_IWL<22510> A_IWL<22509> A_IWL<22508> A_IWL<22507> A_IWL<22506> A_IWL<22505> A_IWL<22504> A_IWL<22503> A_IWL<22502> A_IWL<22501> A_IWL<22500> A_IWL<22499> A_IWL<22498> A_IWL<22497> A_IWL<22496> A_IWL<22495> A_IWL<22494> A_IWL<22493> A_IWL<22492> A_IWL<22491> A_IWL<22490> A_IWL<22489> A_IWL<22488> A_IWL<22487> A_IWL<22486> A_IWL<22485> A_IWL<22484> A_IWL<22483> A_IWL<22482> A_IWL<22481> A_IWL<22480> A_IWL<22479> A_IWL<22478> A_IWL<22477> A_IWL<22476> A_IWL<22475> A_IWL<22474> A_IWL<22473> A_IWL<22472> A_IWL<22471> A_IWL<22470> A_IWL<22469> A_IWL<22468> A_IWL<22467> A_IWL<22466> A_IWL<22465> A_IWL<22464> A_IWL<22463> A_IWL<22462> A_IWL<22461> A_IWL<22460> A_IWL<22459> A_IWL<22458> A_IWL<22457> A_IWL<22456> A_IWL<22455> A_IWL<22454> A_IWL<22453> A_IWL<22452> A_IWL<22451> A_IWL<22450> A_IWL<22449> A_IWL<22448> A_IWL<22447> A_IWL<22446> A_IWL<22445> A_IWL<22444> A_IWL<22443> A_IWL<22442> A_IWL<22441> A_IWL<22440> A_IWL<22439> A_IWL<22438> A_IWL<22437> A_IWL<22436> A_IWL<22435> A_IWL<22434> A_IWL<22433> A_IWL<22432> A_IWL<22431> A_IWL<22430> A_IWL<22429> A_IWL<22428> A_IWL<22427> A_IWL<22426> A_IWL<22425> A_IWL<22424> A_IWL<22423> A_IWL<22422> A_IWL<22421> A_IWL<22420> A_IWL<22419> A_IWL<22418> A_IWL<22417> A_IWL<22416> A_IWL<22415> A_IWL<22414> A_IWL<22413> A_IWL<22412> A_IWL<22411> A_IWL<22410> A_IWL<22409> A_IWL<22408> A_IWL<22407> A_IWL<22406> A_IWL<22405> A_IWL<22404> A_IWL<22403> A_IWL<22402> A_IWL<22401> A_IWL<22400> A_IWL<22399> A_IWL<22398> A_IWL<22397> A_IWL<22396> A_IWL<22395> A_IWL<22394> A_IWL<22393> A_IWL<22392> A_IWL<22391> A_IWL<22390> A_IWL<22389> A_IWL<22388> A_IWL<22387> A_IWL<22386> A_IWL<22385> A_IWL<22384> A_IWL<22383> A_IWL<22382> A_IWL<22381> A_IWL<22380> A_IWL<22379> A_IWL<22378> A_IWL<22377> A_IWL<22376> A_IWL<22375> A_IWL<22374> A_IWL<22373> A_IWL<22372> A_IWL<22371> A_IWL<22370> A_IWL<22369> A_IWL<22368> A_IWL<22367> A_IWL<22366> A_IWL<22365> A_IWL<22364> A_IWL<22363> A_IWL<22362> A_IWL<22361> A_IWL<22360> A_IWL<22359> A_IWL<22358> A_IWL<22357> A_IWL<22356> A_IWL<22355> A_IWL<22354> A_IWL<22353> A_IWL<22352> A_IWL<22351> A_IWL<22350> A_IWL<22349> A_IWL<22348> A_IWL<22347> A_IWL<22346> A_IWL<22345> A_IWL<22344> A_IWL<22343> A_IWL<22342> A_IWL<22341> A_IWL<22340> A_IWL<22339> A_IWL<22338> A_IWL<22337> A_IWL<22336> A_IWL<22335> A_IWL<22334> A_IWL<22333> A_IWL<22332> A_IWL<22331> A_IWL<22330> A_IWL<22329> A_IWL<22328> A_IWL<22327> A_IWL<22326> A_IWL<22325> A_IWL<22324> A_IWL<22323> A_IWL<22322> A_IWL<22321> A_IWL<22320> A_IWL<22319> A_IWL<22318> A_IWL<22317> A_IWL<22316> A_IWL<22315> A_IWL<22314> A_IWL<22313> A_IWL<22312> A_IWL<22311> A_IWL<22310> A_IWL<22309> A_IWL<22308> A_IWL<22307> A_IWL<22306> A_IWL<22305> A_IWL<22304> A_IWL<22303> A_IWL<22302> A_IWL<22301> A_IWL<22300> A_IWL<22299> A_IWL<22298> A_IWL<22297> A_IWL<22296> A_IWL<22295> A_IWL<22294> A_IWL<22293> A_IWL<22292> A_IWL<22291> A_IWL<22290> A_IWL<22289> A_IWL<22288> A_IWL<22287> A_IWL<22286> A_IWL<22285> A_IWL<22284> A_IWL<22283> A_IWL<22282> A_IWL<22281> A_IWL<22280> A_IWL<22279> A_IWL<22278> A_IWL<22277> A_IWL<22276> A_IWL<22275> A_IWL<22274> A_IWL<22273> A_IWL<22272> A_IWL<22271> A_IWL<22270> A_IWL<22269> A_IWL<22268> A_IWL<22267> A_IWL<22266> A_IWL<22265> A_IWL<22264> A_IWL<22263> A_IWL<22262> A_IWL<22261> A_IWL<22260> A_IWL<22259> A_IWL<22258> A_IWL<22257> A_IWL<22256> A_IWL<22255> A_IWL<22254> A_IWL<22253> A_IWL<22252> A_IWL<22251> A_IWL<22250> A_IWL<22249> A_IWL<22248> A_IWL<22247> A_IWL<22246> A_IWL<22245> A_IWL<22244> A_IWL<22243> A_IWL<22242> A_IWL<22241> A_IWL<22240> A_IWL<22239> A_IWL<22238> A_IWL<22237> A_IWL<22236> A_IWL<22235> A_IWL<22234> A_IWL<22233> A_IWL<22232> A_IWL<22231> A_IWL<22230> A_IWL<22229> A_IWL<22228> A_IWL<22227> A_IWL<22226> A_IWL<22225> A_IWL<22224> A_IWL<22223> A_IWL<22222> A_IWL<22221> A_IWL<22220> A_IWL<22219> A_IWL<22218> A_IWL<22217> A_IWL<22216> A_IWL<22215> A_IWL<22214> A_IWL<22213> A_IWL<22212> A_IWL<22211> A_IWL<22210> A_IWL<22209> A_IWL<22208> A_IWL<22207> A_IWL<22206> A_IWL<22205> A_IWL<22204> A_IWL<22203> A_IWL<22202> A_IWL<22201> A_IWL<22200> A_IWL<22199> A_IWL<22198> A_IWL<22197> A_IWL<22196> A_IWL<22195> A_IWL<22194> A_IWL<22193> A_IWL<22192> A_IWL<22191> A_IWL<22190> A_IWL<22189> A_IWL<22188> A_IWL<22187> A_IWL<22186> A_IWL<22185> A_IWL<22184> A_IWL<22183> A_IWL<22182> A_IWL<22181> A_IWL<22180> A_IWL<22179> A_IWL<22178> A_IWL<22177> A_IWL<22176> A_IWL<22175> A_IWL<22174> A_IWL<22173> A_IWL<22172> A_IWL<22171> A_IWL<22170> A_IWL<22169> A_IWL<22168> A_IWL<22167> A_IWL<22166> A_IWL<22165> A_IWL<22164> A_IWL<22163> A_IWL<22162> A_IWL<22161> A_IWL<22160> A_IWL<22159> A_IWL<22158> A_IWL<22157> A_IWL<22156> A_IWL<22155> A_IWL<22154> A_IWL<22153> A_IWL<22152> A_IWL<22151> A_IWL<22150> A_IWL<22149> A_IWL<22148> A_IWL<22147> A_IWL<22146> A_IWL<22145> A_IWL<22144> A_IWL<22143> A_IWL<22142> A_IWL<22141> A_IWL<22140> A_IWL<22139> A_IWL<22138> A_IWL<22137> A_IWL<22136> A_IWL<22135> A_IWL<22134> A_IWL<22133> A_IWL<22132> A_IWL<22131> A_IWL<22130> A_IWL<22129> A_IWL<22128> A_IWL<22127> A_IWL<22126> A_IWL<22125> A_IWL<22124> A_IWL<22123> A_IWL<22122> A_IWL<22121> A_IWL<22120> A_IWL<22119> A_IWL<22118> A_IWL<22117> A_IWL<22116> A_IWL<22115> A_IWL<22114> A_IWL<22113> A_IWL<22112> A_IWL<22111> A_IWL<22110> A_IWL<22109> A_IWL<22108> A_IWL<22107> A_IWL<22106> A_IWL<22105> A_IWL<22104> A_IWL<22103> A_IWL<22102> A_IWL<22101> A_IWL<22100> A_IWL<22099> A_IWL<22098> A_IWL<22097> A_IWL<22096> A_IWL<22095> A_IWL<22094> A_IWL<22093> A_IWL<22092> A_IWL<22091> A_IWL<22090> A_IWL<22089> A_IWL<22088> A_IWL<22087> A_IWL<22086> A_IWL<22085> A_IWL<22084> A_IWL<22083> A_IWL<22082> A_IWL<22081> A_IWL<22080> A_IWL<22079> A_IWL<22078> A_IWL<22077> A_IWL<22076> A_IWL<22075> A_IWL<22074> A_IWL<22073> A_IWL<22072> A_IWL<22071> A_IWL<22070> A_IWL<22069> A_IWL<22068> A_IWL<22067> A_IWL<22066> A_IWL<22065> A_IWL<22064> A_IWL<22063> A_IWL<22062> A_IWL<22061> A_IWL<22060> A_IWL<22059> A_IWL<22058> A_IWL<22057> A_IWL<22056> A_IWL<22055> A_IWL<22054> A_IWL<22053> A_IWL<22052> A_IWL<22051> A_IWL<22050> A_IWL<22049> A_IWL<22048> A_IWL<22047> A_IWL<22046> A_IWL<22045> A_IWL<22044> A_IWL<22043> A_IWL<22042> A_IWL<22041> A_IWL<22040> A_IWL<22039> A_IWL<22038> A_IWL<22037> A_IWL<22036> A_IWL<22035> A_IWL<22034> A_IWL<22033> A_IWL<22032> A_IWL<22031> A_IWL<22030> A_IWL<22029> A_IWL<22028> A_IWL<22027> A_IWL<22026> A_IWL<22025> A_IWL<22024> A_IWL<22023> A_IWL<22022> A_IWL<22021> A_IWL<22020> A_IWL<22019> A_IWL<22018> A_IWL<22017> A_IWL<22016> A_IWL<23039> A_IWL<23038> A_IWL<23037> A_IWL<23036> A_IWL<23035> A_IWL<23034> A_IWL<23033> A_IWL<23032> A_IWL<23031> A_IWL<23030> A_IWL<23029> A_IWL<23028> A_IWL<23027> A_IWL<23026> A_IWL<23025> A_IWL<23024> A_IWL<23023> A_IWL<23022> A_IWL<23021> A_IWL<23020> A_IWL<23019> A_IWL<23018> A_IWL<23017> A_IWL<23016> A_IWL<23015> A_IWL<23014> A_IWL<23013> A_IWL<23012> A_IWL<23011> A_IWL<23010> A_IWL<23009> A_IWL<23008> A_IWL<23007> A_IWL<23006> A_IWL<23005> A_IWL<23004> A_IWL<23003> A_IWL<23002> A_IWL<23001> A_IWL<23000> A_IWL<22999> A_IWL<22998> A_IWL<22997> A_IWL<22996> A_IWL<22995> A_IWL<22994> A_IWL<22993> A_IWL<22992> A_IWL<22991> A_IWL<22990> A_IWL<22989> A_IWL<22988> A_IWL<22987> A_IWL<22986> A_IWL<22985> A_IWL<22984> A_IWL<22983> A_IWL<22982> A_IWL<22981> A_IWL<22980> A_IWL<22979> A_IWL<22978> A_IWL<22977> A_IWL<22976> A_IWL<22975> A_IWL<22974> A_IWL<22973> A_IWL<22972> A_IWL<22971> A_IWL<22970> A_IWL<22969> A_IWL<22968> A_IWL<22967> A_IWL<22966> A_IWL<22965> A_IWL<22964> A_IWL<22963> A_IWL<22962> A_IWL<22961> A_IWL<22960> A_IWL<22959> A_IWL<22958> A_IWL<22957> A_IWL<22956> A_IWL<22955> A_IWL<22954> A_IWL<22953> A_IWL<22952> A_IWL<22951> A_IWL<22950> A_IWL<22949> A_IWL<22948> A_IWL<22947> A_IWL<22946> A_IWL<22945> A_IWL<22944> A_IWL<22943> A_IWL<22942> A_IWL<22941> A_IWL<22940> A_IWL<22939> A_IWL<22938> A_IWL<22937> A_IWL<22936> A_IWL<22935> A_IWL<22934> A_IWL<22933> A_IWL<22932> A_IWL<22931> A_IWL<22930> A_IWL<22929> A_IWL<22928> A_IWL<22927> A_IWL<22926> A_IWL<22925> A_IWL<22924> A_IWL<22923> A_IWL<22922> A_IWL<22921> A_IWL<22920> A_IWL<22919> A_IWL<22918> A_IWL<22917> A_IWL<22916> A_IWL<22915> A_IWL<22914> A_IWL<22913> A_IWL<22912> A_IWL<22911> A_IWL<22910> A_IWL<22909> A_IWL<22908> A_IWL<22907> A_IWL<22906> A_IWL<22905> A_IWL<22904> A_IWL<22903> A_IWL<22902> A_IWL<22901> A_IWL<22900> A_IWL<22899> A_IWL<22898> A_IWL<22897> A_IWL<22896> A_IWL<22895> A_IWL<22894> A_IWL<22893> A_IWL<22892> A_IWL<22891> A_IWL<22890> A_IWL<22889> A_IWL<22888> A_IWL<22887> A_IWL<22886> A_IWL<22885> A_IWL<22884> A_IWL<22883> A_IWL<22882> A_IWL<22881> A_IWL<22880> A_IWL<22879> A_IWL<22878> A_IWL<22877> A_IWL<22876> A_IWL<22875> A_IWL<22874> A_IWL<22873> A_IWL<22872> A_IWL<22871> A_IWL<22870> A_IWL<22869> A_IWL<22868> A_IWL<22867> A_IWL<22866> A_IWL<22865> A_IWL<22864> A_IWL<22863> A_IWL<22862> A_IWL<22861> A_IWL<22860> A_IWL<22859> A_IWL<22858> A_IWL<22857> A_IWL<22856> A_IWL<22855> A_IWL<22854> A_IWL<22853> A_IWL<22852> A_IWL<22851> A_IWL<22850> A_IWL<22849> A_IWL<22848> A_IWL<22847> A_IWL<22846> A_IWL<22845> A_IWL<22844> A_IWL<22843> A_IWL<22842> A_IWL<22841> A_IWL<22840> A_IWL<22839> A_IWL<22838> A_IWL<22837> A_IWL<22836> A_IWL<22835> A_IWL<22834> A_IWL<22833> A_IWL<22832> A_IWL<22831> A_IWL<22830> A_IWL<22829> A_IWL<22828> A_IWL<22827> A_IWL<22826> A_IWL<22825> A_IWL<22824> A_IWL<22823> A_IWL<22822> A_IWL<22821> A_IWL<22820> A_IWL<22819> A_IWL<22818> A_IWL<22817> A_IWL<22816> A_IWL<22815> A_IWL<22814> A_IWL<22813> A_IWL<22812> A_IWL<22811> A_IWL<22810> A_IWL<22809> A_IWL<22808> A_IWL<22807> A_IWL<22806> A_IWL<22805> A_IWL<22804> A_IWL<22803> A_IWL<22802> A_IWL<22801> A_IWL<22800> A_IWL<22799> A_IWL<22798> A_IWL<22797> A_IWL<22796> A_IWL<22795> A_IWL<22794> A_IWL<22793> A_IWL<22792> A_IWL<22791> A_IWL<22790> A_IWL<22789> A_IWL<22788> A_IWL<22787> A_IWL<22786> A_IWL<22785> A_IWL<22784> A_IWL<22783> A_IWL<22782> A_IWL<22781> A_IWL<22780> A_IWL<22779> A_IWL<22778> A_IWL<22777> A_IWL<22776> A_IWL<22775> A_IWL<22774> A_IWL<22773> A_IWL<22772> A_IWL<22771> A_IWL<22770> A_IWL<22769> A_IWL<22768> A_IWL<22767> A_IWL<22766> A_IWL<22765> A_IWL<22764> A_IWL<22763> A_IWL<22762> A_IWL<22761> A_IWL<22760> A_IWL<22759> A_IWL<22758> A_IWL<22757> A_IWL<22756> A_IWL<22755> A_IWL<22754> A_IWL<22753> A_IWL<22752> A_IWL<22751> A_IWL<22750> A_IWL<22749> A_IWL<22748> A_IWL<22747> A_IWL<22746> A_IWL<22745> A_IWL<22744> A_IWL<22743> A_IWL<22742> A_IWL<22741> A_IWL<22740> A_IWL<22739> A_IWL<22738> A_IWL<22737> A_IWL<22736> A_IWL<22735> A_IWL<22734> A_IWL<22733> A_IWL<22732> A_IWL<22731> A_IWL<22730> A_IWL<22729> A_IWL<22728> A_IWL<22727> A_IWL<22726> A_IWL<22725> A_IWL<22724> A_IWL<22723> A_IWL<22722> A_IWL<22721> A_IWL<22720> A_IWL<22719> A_IWL<22718> A_IWL<22717> A_IWL<22716> A_IWL<22715> A_IWL<22714> A_IWL<22713> A_IWL<22712> A_IWL<22711> A_IWL<22710> A_IWL<22709> A_IWL<22708> A_IWL<22707> A_IWL<22706> A_IWL<22705> A_IWL<22704> A_IWL<22703> A_IWL<22702> A_IWL<22701> A_IWL<22700> A_IWL<22699> A_IWL<22698> A_IWL<22697> A_IWL<22696> A_IWL<22695> A_IWL<22694> A_IWL<22693> A_IWL<22692> A_IWL<22691> A_IWL<22690> A_IWL<22689> A_IWL<22688> A_IWL<22687> A_IWL<22686> A_IWL<22685> A_IWL<22684> A_IWL<22683> A_IWL<22682> A_IWL<22681> A_IWL<22680> A_IWL<22679> A_IWL<22678> A_IWL<22677> A_IWL<22676> A_IWL<22675> A_IWL<22674> A_IWL<22673> A_IWL<22672> A_IWL<22671> A_IWL<22670> A_IWL<22669> A_IWL<22668> A_IWL<22667> A_IWL<22666> A_IWL<22665> A_IWL<22664> A_IWL<22663> A_IWL<22662> A_IWL<22661> A_IWL<22660> A_IWL<22659> A_IWL<22658> A_IWL<22657> A_IWL<22656> A_IWL<22655> A_IWL<22654> A_IWL<22653> A_IWL<22652> A_IWL<22651> A_IWL<22650> A_IWL<22649> A_IWL<22648> A_IWL<22647> A_IWL<22646> A_IWL<22645> A_IWL<22644> A_IWL<22643> A_IWL<22642> A_IWL<22641> A_IWL<22640> A_IWL<22639> A_IWL<22638> A_IWL<22637> A_IWL<22636> A_IWL<22635> A_IWL<22634> A_IWL<22633> A_IWL<22632> A_IWL<22631> A_IWL<22630> A_IWL<22629> A_IWL<22628> A_IWL<22627> A_IWL<22626> A_IWL<22625> A_IWL<22624> A_IWL<22623> A_IWL<22622> A_IWL<22621> A_IWL<22620> A_IWL<22619> A_IWL<22618> A_IWL<22617> A_IWL<22616> A_IWL<22615> A_IWL<22614> A_IWL<22613> A_IWL<22612> A_IWL<22611> A_IWL<22610> A_IWL<22609> A_IWL<22608> A_IWL<22607> A_IWL<22606> A_IWL<22605> A_IWL<22604> A_IWL<22603> A_IWL<22602> A_IWL<22601> A_IWL<22600> A_IWL<22599> A_IWL<22598> A_IWL<22597> A_IWL<22596> A_IWL<22595> A_IWL<22594> A_IWL<22593> A_IWL<22592> A_IWL<22591> A_IWL<22590> A_IWL<22589> A_IWL<22588> A_IWL<22587> A_IWL<22586> A_IWL<22585> A_IWL<22584> A_IWL<22583> A_IWL<22582> A_IWL<22581> A_IWL<22580> A_IWL<22579> A_IWL<22578> A_IWL<22577> A_IWL<22576> A_IWL<22575> A_IWL<22574> A_IWL<22573> A_IWL<22572> A_IWL<22571> A_IWL<22570> A_IWL<22569> A_IWL<22568> A_IWL<22567> A_IWL<22566> A_IWL<22565> A_IWL<22564> A_IWL<22563> A_IWL<22562> A_IWL<22561> A_IWL<22560> A_IWL<22559> A_IWL<22558> A_IWL<22557> A_IWL<22556> A_IWL<22555> A_IWL<22554> A_IWL<22553> A_IWL<22552> A_IWL<22551> A_IWL<22550> A_IWL<22549> A_IWL<22548> A_IWL<22547> A_IWL<22546> A_IWL<22545> A_IWL<22544> A_IWL<22543> A_IWL<22542> A_IWL<22541> A_IWL<22540> A_IWL<22539> A_IWL<22538> A_IWL<22537> A_IWL<22536> A_IWL<22535> A_IWL<22534> A_IWL<22533> A_IWL<22532> A_IWL<22531> A_IWL<22530> A_IWL<22529> A_IWL<22528> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<43> A_BLC<87> A_BLC<86> A_BLC_TOP<87> A_BLC_TOP<86> A_BLT<87> A_BLT<86> A_BLT_TOP<87> A_BLT_TOP<86> A_IWL<22015> A_IWL<22014> A_IWL<22013> A_IWL<22012> A_IWL<22011> A_IWL<22010> A_IWL<22009> A_IWL<22008> A_IWL<22007> A_IWL<22006> A_IWL<22005> A_IWL<22004> A_IWL<22003> A_IWL<22002> A_IWL<22001> A_IWL<22000> A_IWL<21999> A_IWL<21998> A_IWL<21997> A_IWL<21996> A_IWL<21995> A_IWL<21994> A_IWL<21993> A_IWL<21992> A_IWL<21991> A_IWL<21990> A_IWL<21989> A_IWL<21988> A_IWL<21987> A_IWL<21986> A_IWL<21985> A_IWL<21984> A_IWL<21983> A_IWL<21982> A_IWL<21981> A_IWL<21980> A_IWL<21979> A_IWL<21978> A_IWL<21977> A_IWL<21976> A_IWL<21975> A_IWL<21974> A_IWL<21973> A_IWL<21972> A_IWL<21971> A_IWL<21970> A_IWL<21969> A_IWL<21968> A_IWL<21967> A_IWL<21966> A_IWL<21965> A_IWL<21964> A_IWL<21963> A_IWL<21962> A_IWL<21961> A_IWL<21960> A_IWL<21959> A_IWL<21958> A_IWL<21957> A_IWL<21956> A_IWL<21955> A_IWL<21954> A_IWL<21953> A_IWL<21952> A_IWL<21951> A_IWL<21950> A_IWL<21949> A_IWL<21948> A_IWL<21947> A_IWL<21946> A_IWL<21945> A_IWL<21944> A_IWL<21943> A_IWL<21942> A_IWL<21941> A_IWL<21940> A_IWL<21939> A_IWL<21938> A_IWL<21937> A_IWL<21936> A_IWL<21935> A_IWL<21934> A_IWL<21933> A_IWL<21932> A_IWL<21931> A_IWL<21930> A_IWL<21929> A_IWL<21928> A_IWL<21927> A_IWL<21926> A_IWL<21925> A_IWL<21924> A_IWL<21923> A_IWL<21922> A_IWL<21921> A_IWL<21920> A_IWL<21919> A_IWL<21918> A_IWL<21917> A_IWL<21916> A_IWL<21915> A_IWL<21914> A_IWL<21913> A_IWL<21912> A_IWL<21911> A_IWL<21910> A_IWL<21909> A_IWL<21908> A_IWL<21907> A_IWL<21906> A_IWL<21905> A_IWL<21904> A_IWL<21903> A_IWL<21902> A_IWL<21901> A_IWL<21900> A_IWL<21899> A_IWL<21898> A_IWL<21897> A_IWL<21896> A_IWL<21895> A_IWL<21894> A_IWL<21893> A_IWL<21892> A_IWL<21891> A_IWL<21890> A_IWL<21889> A_IWL<21888> A_IWL<21887> A_IWL<21886> A_IWL<21885> A_IWL<21884> A_IWL<21883> A_IWL<21882> A_IWL<21881> A_IWL<21880> A_IWL<21879> A_IWL<21878> A_IWL<21877> A_IWL<21876> A_IWL<21875> A_IWL<21874> A_IWL<21873> A_IWL<21872> A_IWL<21871> A_IWL<21870> A_IWL<21869> A_IWL<21868> A_IWL<21867> A_IWL<21866> A_IWL<21865> A_IWL<21864> A_IWL<21863> A_IWL<21862> A_IWL<21861> A_IWL<21860> A_IWL<21859> A_IWL<21858> A_IWL<21857> A_IWL<21856> A_IWL<21855> A_IWL<21854> A_IWL<21853> A_IWL<21852> A_IWL<21851> A_IWL<21850> A_IWL<21849> A_IWL<21848> A_IWL<21847> A_IWL<21846> A_IWL<21845> A_IWL<21844> A_IWL<21843> A_IWL<21842> A_IWL<21841> A_IWL<21840> A_IWL<21839> A_IWL<21838> A_IWL<21837> A_IWL<21836> A_IWL<21835> A_IWL<21834> A_IWL<21833> A_IWL<21832> A_IWL<21831> A_IWL<21830> A_IWL<21829> A_IWL<21828> A_IWL<21827> A_IWL<21826> A_IWL<21825> A_IWL<21824> A_IWL<21823> A_IWL<21822> A_IWL<21821> A_IWL<21820> A_IWL<21819> A_IWL<21818> A_IWL<21817> A_IWL<21816> A_IWL<21815> A_IWL<21814> A_IWL<21813> A_IWL<21812> A_IWL<21811> A_IWL<21810> A_IWL<21809> A_IWL<21808> A_IWL<21807> A_IWL<21806> A_IWL<21805> A_IWL<21804> A_IWL<21803> A_IWL<21802> A_IWL<21801> A_IWL<21800> A_IWL<21799> A_IWL<21798> A_IWL<21797> A_IWL<21796> A_IWL<21795> A_IWL<21794> A_IWL<21793> A_IWL<21792> A_IWL<21791> A_IWL<21790> A_IWL<21789> A_IWL<21788> A_IWL<21787> A_IWL<21786> A_IWL<21785> A_IWL<21784> A_IWL<21783> A_IWL<21782> A_IWL<21781> A_IWL<21780> A_IWL<21779> A_IWL<21778> A_IWL<21777> A_IWL<21776> A_IWL<21775> A_IWL<21774> A_IWL<21773> A_IWL<21772> A_IWL<21771> A_IWL<21770> A_IWL<21769> A_IWL<21768> A_IWL<21767> A_IWL<21766> A_IWL<21765> A_IWL<21764> A_IWL<21763> A_IWL<21762> A_IWL<21761> A_IWL<21760> A_IWL<21759> A_IWL<21758> A_IWL<21757> A_IWL<21756> A_IWL<21755> A_IWL<21754> A_IWL<21753> A_IWL<21752> A_IWL<21751> A_IWL<21750> A_IWL<21749> A_IWL<21748> A_IWL<21747> A_IWL<21746> A_IWL<21745> A_IWL<21744> A_IWL<21743> A_IWL<21742> A_IWL<21741> A_IWL<21740> A_IWL<21739> A_IWL<21738> A_IWL<21737> A_IWL<21736> A_IWL<21735> A_IWL<21734> A_IWL<21733> A_IWL<21732> A_IWL<21731> A_IWL<21730> A_IWL<21729> A_IWL<21728> A_IWL<21727> A_IWL<21726> A_IWL<21725> A_IWL<21724> A_IWL<21723> A_IWL<21722> A_IWL<21721> A_IWL<21720> A_IWL<21719> A_IWL<21718> A_IWL<21717> A_IWL<21716> A_IWL<21715> A_IWL<21714> A_IWL<21713> A_IWL<21712> A_IWL<21711> A_IWL<21710> A_IWL<21709> A_IWL<21708> A_IWL<21707> A_IWL<21706> A_IWL<21705> A_IWL<21704> A_IWL<21703> A_IWL<21702> A_IWL<21701> A_IWL<21700> A_IWL<21699> A_IWL<21698> A_IWL<21697> A_IWL<21696> A_IWL<21695> A_IWL<21694> A_IWL<21693> A_IWL<21692> A_IWL<21691> A_IWL<21690> A_IWL<21689> A_IWL<21688> A_IWL<21687> A_IWL<21686> A_IWL<21685> A_IWL<21684> A_IWL<21683> A_IWL<21682> A_IWL<21681> A_IWL<21680> A_IWL<21679> A_IWL<21678> A_IWL<21677> A_IWL<21676> A_IWL<21675> A_IWL<21674> A_IWL<21673> A_IWL<21672> A_IWL<21671> A_IWL<21670> A_IWL<21669> A_IWL<21668> A_IWL<21667> A_IWL<21666> A_IWL<21665> A_IWL<21664> A_IWL<21663> A_IWL<21662> A_IWL<21661> A_IWL<21660> A_IWL<21659> A_IWL<21658> A_IWL<21657> A_IWL<21656> A_IWL<21655> A_IWL<21654> A_IWL<21653> A_IWL<21652> A_IWL<21651> A_IWL<21650> A_IWL<21649> A_IWL<21648> A_IWL<21647> A_IWL<21646> A_IWL<21645> A_IWL<21644> A_IWL<21643> A_IWL<21642> A_IWL<21641> A_IWL<21640> A_IWL<21639> A_IWL<21638> A_IWL<21637> A_IWL<21636> A_IWL<21635> A_IWL<21634> A_IWL<21633> A_IWL<21632> A_IWL<21631> A_IWL<21630> A_IWL<21629> A_IWL<21628> A_IWL<21627> A_IWL<21626> A_IWL<21625> A_IWL<21624> A_IWL<21623> A_IWL<21622> A_IWL<21621> A_IWL<21620> A_IWL<21619> A_IWL<21618> A_IWL<21617> A_IWL<21616> A_IWL<21615> A_IWL<21614> A_IWL<21613> A_IWL<21612> A_IWL<21611> A_IWL<21610> A_IWL<21609> A_IWL<21608> A_IWL<21607> A_IWL<21606> A_IWL<21605> A_IWL<21604> A_IWL<21603> A_IWL<21602> A_IWL<21601> A_IWL<21600> A_IWL<21599> A_IWL<21598> A_IWL<21597> A_IWL<21596> A_IWL<21595> A_IWL<21594> A_IWL<21593> A_IWL<21592> A_IWL<21591> A_IWL<21590> A_IWL<21589> A_IWL<21588> A_IWL<21587> A_IWL<21586> A_IWL<21585> A_IWL<21584> A_IWL<21583> A_IWL<21582> A_IWL<21581> A_IWL<21580> A_IWL<21579> A_IWL<21578> A_IWL<21577> A_IWL<21576> A_IWL<21575> A_IWL<21574> A_IWL<21573> A_IWL<21572> A_IWL<21571> A_IWL<21570> A_IWL<21569> A_IWL<21568> A_IWL<21567> A_IWL<21566> A_IWL<21565> A_IWL<21564> A_IWL<21563> A_IWL<21562> A_IWL<21561> A_IWL<21560> A_IWL<21559> A_IWL<21558> A_IWL<21557> A_IWL<21556> A_IWL<21555> A_IWL<21554> A_IWL<21553> A_IWL<21552> A_IWL<21551> A_IWL<21550> A_IWL<21549> A_IWL<21548> A_IWL<21547> A_IWL<21546> A_IWL<21545> A_IWL<21544> A_IWL<21543> A_IWL<21542> A_IWL<21541> A_IWL<21540> A_IWL<21539> A_IWL<21538> A_IWL<21537> A_IWL<21536> A_IWL<21535> A_IWL<21534> A_IWL<21533> A_IWL<21532> A_IWL<21531> A_IWL<21530> A_IWL<21529> A_IWL<21528> A_IWL<21527> A_IWL<21526> A_IWL<21525> A_IWL<21524> A_IWL<21523> A_IWL<21522> A_IWL<21521> A_IWL<21520> A_IWL<21519> A_IWL<21518> A_IWL<21517> A_IWL<21516> A_IWL<21515> A_IWL<21514> A_IWL<21513> A_IWL<21512> A_IWL<21511> A_IWL<21510> A_IWL<21509> A_IWL<21508> A_IWL<21507> A_IWL<21506> A_IWL<21505> A_IWL<21504> A_IWL<22527> A_IWL<22526> A_IWL<22525> A_IWL<22524> A_IWL<22523> A_IWL<22522> A_IWL<22521> A_IWL<22520> A_IWL<22519> A_IWL<22518> A_IWL<22517> A_IWL<22516> A_IWL<22515> A_IWL<22514> A_IWL<22513> A_IWL<22512> A_IWL<22511> A_IWL<22510> A_IWL<22509> A_IWL<22508> A_IWL<22507> A_IWL<22506> A_IWL<22505> A_IWL<22504> A_IWL<22503> A_IWL<22502> A_IWL<22501> A_IWL<22500> A_IWL<22499> A_IWL<22498> A_IWL<22497> A_IWL<22496> A_IWL<22495> A_IWL<22494> A_IWL<22493> A_IWL<22492> A_IWL<22491> A_IWL<22490> A_IWL<22489> A_IWL<22488> A_IWL<22487> A_IWL<22486> A_IWL<22485> A_IWL<22484> A_IWL<22483> A_IWL<22482> A_IWL<22481> A_IWL<22480> A_IWL<22479> A_IWL<22478> A_IWL<22477> A_IWL<22476> A_IWL<22475> A_IWL<22474> A_IWL<22473> A_IWL<22472> A_IWL<22471> A_IWL<22470> A_IWL<22469> A_IWL<22468> A_IWL<22467> A_IWL<22466> A_IWL<22465> A_IWL<22464> A_IWL<22463> A_IWL<22462> A_IWL<22461> A_IWL<22460> A_IWL<22459> A_IWL<22458> A_IWL<22457> A_IWL<22456> A_IWL<22455> A_IWL<22454> A_IWL<22453> A_IWL<22452> A_IWL<22451> A_IWL<22450> A_IWL<22449> A_IWL<22448> A_IWL<22447> A_IWL<22446> A_IWL<22445> A_IWL<22444> A_IWL<22443> A_IWL<22442> A_IWL<22441> A_IWL<22440> A_IWL<22439> A_IWL<22438> A_IWL<22437> A_IWL<22436> A_IWL<22435> A_IWL<22434> A_IWL<22433> A_IWL<22432> A_IWL<22431> A_IWL<22430> A_IWL<22429> A_IWL<22428> A_IWL<22427> A_IWL<22426> A_IWL<22425> A_IWL<22424> A_IWL<22423> A_IWL<22422> A_IWL<22421> A_IWL<22420> A_IWL<22419> A_IWL<22418> A_IWL<22417> A_IWL<22416> A_IWL<22415> A_IWL<22414> A_IWL<22413> A_IWL<22412> A_IWL<22411> A_IWL<22410> A_IWL<22409> A_IWL<22408> A_IWL<22407> A_IWL<22406> A_IWL<22405> A_IWL<22404> A_IWL<22403> A_IWL<22402> A_IWL<22401> A_IWL<22400> A_IWL<22399> A_IWL<22398> A_IWL<22397> A_IWL<22396> A_IWL<22395> A_IWL<22394> A_IWL<22393> A_IWL<22392> A_IWL<22391> A_IWL<22390> A_IWL<22389> A_IWL<22388> A_IWL<22387> A_IWL<22386> A_IWL<22385> A_IWL<22384> A_IWL<22383> A_IWL<22382> A_IWL<22381> A_IWL<22380> A_IWL<22379> A_IWL<22378> A_IWL<22377> A_IWL<22376> A_IWL<22375> A_IWL<22374> A_IWL<22373> A_IWL<22372> A_IWL<22371> A_IWL<22370> A_IWL<22369> A_IWL<22368> A_IWL<22367> A_IWL<22366> A_IWL<22365> A_IWL<22364> A_IWL<22363> A_IWL<22362> A_IWL<22361> A_IWL<22360> A_IWL<22359> A_IWL<22358> A_IWL<22357> A_IWL<22356> A_IWL<22355> A_IWL<22354> A_IWL<22353> A_IWL<22352> A_IWL<22351> A_IWL<22350> A_IWL<22349> A_IWL<22348> A_IWL<22347> A_IWL<22346> A_IWL<22345> A_IWL<22344> A_IWL<22343> A_IWL<22342> A_IWL<22341> A_IWL<22340> A_IWL<22339> A_IWL<22338> A_IWL<22337> A_IWL<22336> A_IWL<22335> A_IWL<22334> A_IWL<22333> A_IWL<22332> A_IWL<22331> A_IWL<22330> A_IWL<22329> A_IWL<22328> A_IWL<22327> A_IWL<22326> A_IWL<22325> A_IWL<22324> A_IWL<22323> A_IWL<22322> A_IWL<22321> A_IWL<22320> A_IWL<22319> A_IWL<22318> A_IWL<22317> A_IWL<22316> A_IWL<22315> A_IWL<22314> A_IWL<22313> A_IWL<22312> A_IWL<22311> A_IWL<22310> A_IWL<22309> A_IWL<22308> A_IWL<22307> A_IWL<22306> A_IWL<22305> A_IWL<22304> A_IWL<22303> A_IWL<22302> A_IWL<22301> A_IWL<22300> A_IWL<22299> A_IWL<22298> A_IWL<22297> A_IWL<22296> A_IWL<22295> A_IWL<22294> A_IWL<22293> A_IWL<22292> A_IWL<22291> A_IWL<22290> A_IWL<22289> A_IWL<22288> A_IWL<22287> A_IWL<22286> A_IWL<22285> A_IWL<22284> A_IWL<22283> A_IWL<22282> A_IWL<22281> A_IWL<22280> A_IWL<22279> A_IWL<22278> A_IWL<22277> A_IWL<22276> A_IWL<22275> A_IWL<22274> A_IWL<22273> A_IWL<22272> A_IWL<22271> A_IWL<22270> A_IWL<22269> A_IWL<22268> A_IWL<22267> A_IWL<22266> A_IWL<22265> A_IWL<22264> A_IWL<22263> A_IWL<22262> A_IWL<22261> A_IWL<22260> A_IWL<22259> A_IWL<22258> A_IWL<22257> A_IWL<22256> A_IWL<22255> A_IWL<22254> A_IWL<22253> A_IWL<22252> A_IWL<22251> A_IWL<22250> A_IWL<22249> A_IWL<22248> A_IWL<22247> A_IWL<22246> A_IWL<22245> A_IWL<22244> A_IWL<22243> A_IWL<22242> A_IWL<22241> A_IWL<22240> A_IWL<22239> A_IWL<22238> A_IWL<22237> A_IWL<22236> A_IWL<22235> A_IWL<22234> A_IWL<22233> A_IWL<22232> A_IWL<22231> A_IWL<22230> A_IWL<22229> A_IWL<22228> A_IWL<22227> A_IWL<22226> A_IWL<22225> A_IWL<22224> A_IWL<22223> A_IWL<22222> A_IWL<22221> A_IWL<22220> A_IWL<22219> A_IWL<22218> A_IWL<22217> A_IWL<22216> A_IWL<22215> A_IWL<22214> A_IWL<22213> A_IWL<22212> A_IWL<22211> A_IWL<22210> A_IWL<22209> A_IWL<22208> A_IWL<22207> A_IWL<22206> A_IWL<22205> A_IWL<22204> A_IWL<22203> A_IWL<22202> A_IWL<22201> A_IWL<22200> A_IWL<22199> A_IWL<22198> A_IWL<22197> A_IWL<22196> A_IWL<22195> A_IWL<22194> A_IWL<22193> A_IWL<22192> A_IWL<22191> A_IWL<22190> A_IWL<22189> A_IWL<22188> A_IWL<22187> A_IWL<22186> A_IWL<22185> A_IWL<22184> A_IWL<22183> A_IWL<22182> A_IWL<22181> A_IWL<22180> A_IWL<22179> A_IWL<22178> A_IWL<22177> A_IWL<22176> A_IWL<22175> A_IWL<22174> A_IWL<22173> A_IWL<22172> A_IWL<22171> A_IWL<22170> A_IWL<22169> A_IWL<22168> A_IWL<22167> A_IWL<22166> A_IWL<22165> A_IWL<22164> A_IWL<22163> A_IWL<22162> A_IWL<22161> A_IWL<22160> A_IWL<22159> A_IWL<22158> A_IWL<22157> A_IWL<22156> A_IWL<22155> A_IWL<22154> A_IWL<22153> A_IWL<22152> A_IWL<22151> A_IWL<22150> A_IWL<22149> A_IWL<22148> A_IWL<22147> A_IWL<22146> A_IWL<22145> A_IWL<22144> A_IWL<22143> A_IWL<22142> A_IWL<22141> A_IWL<22140> A_IWL<22139> A_IWL<22138> A_IWL<22137> A_IWL<22136> A_IWL<22135> A_IWL<22134> A_IWL<22133> A_IWL<22132> A_IWL<22131> A_IWL<22130> A_IWL<22129> A_IWL<22128> A_IWL<22127> A_IWL<22126> A_IWL<22125> A_IWL<22124> A_IWL<22123> A_IWL<22122> A_IWL<22121> A_IWL<22120> A_IWL<22119> A_IWL<22118> A_IWL<22117> A_IWL<22116> A_IWL<22115> A_IWL<22114> A_IWL<22113> A_IWL<22112> A_IWL<22111> A_IWL<22110> A_IWL<22109> A_IWL<22108> A_IWL<22107> A_IWL<22106> A_IWL<22105> A_IWL<22104> A_IWL<22103> A_IWL<22102> A_IWL<22101> A_IWL<22100> A_IWL<22099> A_IWL<22098> A_IWL<22097> A_IWL<22096> A_IWL<22095> A_IWL<22094> A_IWL<22093> A_IWL<22092> A_IWL<22091> A_IWL<22090> A_IWL<22089> A_IWL<22088> A_IWL<22087> A_IWL<22086> A_IWL<22085> A_IWL<22084> A_IWL<22083> A_IWL<22082> A_IWL<22081> A_IWL<22080> A_IWL<22079> A_IWL<22078> A_IWL<22077> A_IWL<22076> A_IWL<22075> A_IWL<22074> A_IWL<22073> A_IWL<22072> A_IWL<22071> A_IWL<22070> A_IWL<22069> A_IWL<22068> A_IWL<22067> A_IWL<22066> A_IWL<22065> A_IWL<22064> A_IWL<22063> A_IWL<22062> A_IWL<22061> A_IWL<22060> A_IWL<22059> A_IWL<22058> A_IWL<22057> A_IWL<22056> A_IWL<22055> A_IWL<22054> A_IWL<22053> A_IWL<22052> A_IWL<22051> A_IWL<22050> A_IWL<22049> A_IWL<22048> A_IWL<22047> A_IWL<22046> A_IWL<22045> A_IWL<22044> A_IWL<22043> A_IWL<22042> A_IWL<22041> A_IWL<22040> A_IWL<22039> A_IWL<22038> A_IWL<22037> A_IWL<22036> A_IWL<22035> A_IWL<22034> A_IWL<22033> A_IWL<22032> A_IWL<22031> A_IWL<22030> A_IWL<22029> A_IWL<22028> A_IWL<22027> A_IWL<22026> A_IWL<22025> A_IWL<22024> A_IWL<22023> A_IWL<22022> A_IWL<22021> A_IWL<22020> A_IWL<22019> A_IWL<22018> A_IWL<22017> A_IWL<22016> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<42> A_BLC<85> A_BLC<84> A_BLC_TOP<85> A_BLC_TOP<84> A_BLT<85> A_BLT<84> A_BLT_TOP<85> A_BLT_TOP<84> A_IWL<21503> A_IWL<21502> A_IWL<21501> A_IWL<21500> A_IWL<21499> A_IWL<21498> A_IWL<21497> A_IWL<21496> A_IWL<21495> A_IWL<21494> A_IWL<21493> A_IWL<21492> A_IWL<21491> A_IWL<21490> A_IWL<21489> A_IWL<21488> A_IWL<21487> A_IWL<21486> A_IWL<21485> A_IWL<21484> A_IWL<21483> A_IWL<21482> A_IWL<21481> A_IWL<21480> A_IWL<21479> A_IWL<21478> A_IWL<21477> A_IWL<21476> A_IWL<21475> A_IWL<21474> A_IWL<21473> A_IWL<21472> A_IWL<21471> A_IWL<21470> A_IWL<21469> A_IWL<21468> A_IWL<21467> A_IWL<21466> A_IWL<21465> A_IWL<21464> A_IWL<21463> A_IWL<21462> A_IWL<21461> A_IWL<21460> A_IWL<21459> A_IWL<21458> A_IWL<21457> A_IWL<21456> A_IWL<21455> A_IWL<21454> A_IWL<21453> A_IWL<21452> A_IWL<21451> A_IWL<21450> A_IWL<21449> A_IWL<21448> A_IWL<21447> A_IWL<21446> A_IWL<21445> A_IWL<21444> A_IWL<21443> A_IWL<21442> A_IWL<21441> A_IWL<21440> A_IWL<21439> A_IWL<21438> A_IWL<21437> A_IWL<21436> A_IWL<21435> A_IWL<21434> A_IWL<21433> A_IWL<21432> A_IWL<21431> A_IWL<21430> A_IWL<21429> A_IWL<21428> A_IWL<21427> A_IWL<21426> A_IWL<21425> A_IWL<21424> A_IWL<21423> A_IWL<21422> A_IWL<21421> A_IWL<21420> A_IWL<21419> A_IWL<21418> A_IWL<21417> A_IWL<21416> A_IWL<21415> A_IWL<21414> A_IWL<21413> A_IWL<21412> A_IWL<21411> A_IWL<21410> A_IWL<21409> A_IWL<21408> A_IWL<21407> A_IWL<21406> A_IWL<21405> A_IWL<21404> A_IWL<21403> A_IWL<21402> A_IWL<21401> A_IWL<21400> A_IWL<21399> A_IWL<21398> A_IWL<21397> A_IWL<21396> A_IWL<21395> A_IWL<21394> A_IWL<21393> A_IWL<21392> A_IWL<21391> A_IWL<21390> A_IWL<21389> A_IWL<21388> A_IWL<21387> A_IWL<21386> A_IWL<21385> A_IWL<21384> A_IWL<21383> A_IWL<21382> A_IWL<21381> A_IWL<21380> A_IWL<21379> A_IWL<21378> A_IWL<21377> A_IWL<21376> A_IWL<21375> A_IWL<21374> A_IWL<21373> A_IWL<21372> A_IWL<21371> A_IWL<21370> A_IWL<21369> A_IWL<21368> A_IWL<21367> A_IWL<21366> A_IWL<21365> A_IWL<21364> A_IWL<21363> A_IWL<21362> A_IWL<21361> A_IWL<21360> A_IWL<21359> A_IWL<21358> A_IWL<21357> A_IWL<21356> A_IWL<21355> A_IWL<21354> A_IWL<21353> A_IWL<21352> A_IWL<21351> A_IWL<21350> A_IWL<21349> A_IWL<21348> A_IWL<21347> A_IWL<21346> A_IWL<21345> A_IWL<21344> A_IWL<21343> A_IWL<21342> A_IWL<21341> A_IWL<21340> A_IWL<21339> A_IWL<21338> A_IWL<21337> A_IWL<21336> A_IWL<21335> A_IWL<21334> A_IWL<21333> A_IWL<21332> A_IWL<21331> A_IWL<21330> A_IWL<21329> A_IWL<21328> A_IWL<21327> A_IWL<21326> A_IWL<21325> A_IWL<21324> A_IWL<21323> A_IWL<21322> A_IWL<21321> A_IWL<21320> A_IWL<21319> A_IWL<21318> A_IWL<21317> A_IWL<21316> A_IWL<21315> A_IWL<21314> A_IWL<21313> A_IWL<21312> A_IWL<21311> A_IWL<21310> A_IWL<21309> A_IWL<21308> A_IWL<21307> A_IWL<21306> A_IWL<21305> A_IWL<21304> A_IWL<21303> A_IWL<21302> A_IWL<21301> A_IWL<21300> A_IWL<21299> A_IWL<21298> A_IWL<21297> A_IWL<21296> A_IWL<21295> A_IWL<21294> A_IWL<21293> A_IWL<21292> A_IWL<21291> A_IWL<21290> A_IWL<21289> A_IWL<21288> A_IWL<21287> A_IWL<21286> A_IWL<21285> A_IWL<21284> A_IWL<21283> A_IWL<21282> A_IWL<21281> A_IWL<21280> A_IWL<21279> A_IWL<21278> A_IWL<21277> A_IWL<21276> A_IWL<21275> A_IWL<21274> A_IWL<21273> A_IWL<21272> A_IWL<21271> A_IWL<21270> A_IWL<21269> A_IWL<21268> A_IWL<21267> A_IWL<21266> A_IWL<21265> A_IWL<21264> A_IWL<21263> A_IWL<21262> A_IWL<21261> A_IWL<21260> A_IWL<21259> A_IWL<21258> A_IWL<21257> A_IWL<21256> A_IWL<21255> A_IWL<21254> A_IWL<21253> A_IWL<21252> A_IWL<21251> A_IWL<21250> A_IWL<21249> A_IWL<21248> A_IWL<21247> A_IWL<21246> A_IWL<21245> A_IWL<21244> A_IWL<21243> A_IWL<21242> A_IWL<21241> A_IWL<21240> A_IWL<21239> A_IWL<21238> A_IWL<21237> A_IWL<21236> A_IWL<21235> A_IWL<21234> A_IWL<21233> A_IWL<21232> A_IWL<21231> A_IWL<21230> A_IWL<21229> A_IWL<21228> A_IWL<21227> A_IWL<21226> A_IWL<21225> A_IWL<21224> A_IWL<21223> A_IWL<21222> A_IWL<21221> A_IWL<21220> A_IWL<21219> A_IWL<21218> A_IWL<21217> A_IWL<21216> A_IWL<21215> A_IWL<21214> A_IWL<21213> A_IWL<21212> A_IWL<21211> A_IWL<21210> A_IWL<21209> A_IWL<21208> A_IWL<21207> A_IWL<21206> A_IWL<21205> A_IWL<21204> A_IWL<21203> A_IWL<21202> A_IWL<21201> A_IWL<21200> A_IWL<21199> A_IWL<21198> A_IWL<21197> A_IWL<21196> A_IWL<21195> A_IWL<21194> A_IWL<21193> A_IWL<21192> A_IWL<21191> A_IWL<21190> A_IWL<21189> A_IWL<21188> A_IWL<21187> A_IWL<21186> A_IWL<21185> A_IWL<21184> A_IWL<21183> A_IWL<21182> A_IWL<21181> A_IWL<21180> A_IWL<21179> A_IWL<21178> A_IWL<21177> A_IWL<21176> A_IWL<21175> A_IWL<21174> A_IWL<21173> A_IWL<21172> A_IWL<21171> A_IWL<21170> A_IWL<21169> A_IWL<21168> A_IWL<21167> A_IWL<21166> A_IWL<21165> A_IWL<21164> A_IWL<21163> A_IWL<21162> A_IWL<21161> A_IWL<21160> A_IWL<21159> A_IWL<21158> A_IWL<21157> A_IWL<21156> A_IWL<21155> A_IWL<21154> A_IWL<21153> A_IWL<21152> A_IWL<21151> A_IWL<21150> A_IWL<21149> A_IWL<21148> A_IWL<21147> A_IWL<21146> A_IWL<21145> A_IWL<21144> A_IWL<21143> A_IWL<21142> A_IWL<21141> A_IWL<21140> A_IWL<21139> A_IWL<21138> A_IWL<21137> A_IWL<21136> A_IWL<21135> A_IWL<21134> A_IWL<21133> A_IWL<21132> A_IWL<21131> A_IWL<21130> A_IWL<21129> A_IWL<21128> A_IWL<21127> A_IWL<21126> A_IWL<21125> A_IWL<21124> A_IWL<21123> A_IWL<21122> A_IWL<21121> A_IWL<21120> A_IWL<21119> A_IWL<21118> A_IWL<21117> A_IWL<21116> A_IWL<21115> A_IWL<21114> A_IWL<21113> A_IWL<21112> A_IWL<21111> A_IWL<21110> A_IWL<21109> A_IWL<21108> A_IWL<21107> A_IWL<21106> A_IWL<21105> A_IWL<21104> A_IWL<21103> A_IWL<21102> A_IWL<21101> A_IWL<21100> A_IWL<21099> A_IWL<21098> A_IWL<21097> A_IWL<21096> A_IWL<21095> A_IWL<21094> A_IWL<21093> A_IWL<21092> A_IWL<21091> A_IWL<21090> A_IWL<21089> A_IWL<21088> A_IWL<21087> A_IWL<21086> A_IWL<21085> A_IWL<21084> A_IWL<21083> A_IWL<21082> A_IWL<21081> A_IWL<21080> A_IWL<21079> A_IWL<21078> A_IWL<21077> A_IWL<21076> A_IWL<21075> A_IWL<21074> A_IWL<21073> A_IWL<21072> A_IWL<21071> A_IWL<21070> A_IWL<21069> A_IWL<21068> A_IWL<21067> A_IWL<21066> A_IWL<21065> A_IWL<21064> A_IWL<21063> A_IWL<21062> A_IWL<21061> A_IWL<21060> A_IWL<21059> A_IWL<21058> A_IWL<21057> A_IWL<21056> A_IWL<21055> A_IWL<21054> A_IWL<21053> A_IWL<21052> A_IWL<21051> A_IWL<21050> A_IWL<21049> A_IWL<21048> A_IWL<21047> A_IWL<21046> A_IWL<21045> A_IWL<21044> A_IWL<21043> A_IWL<21042> A_IWL<21041> A_IWL<21040> A_IWL<21039> A_IWL<21038> A_IWL<21037> A_IWL<21036> A_IWL<21035> A_IWL<21034> A_IWL<21033> A_IWL<21032> A_IWL<21031> A_IWL<21030> A_IWL<21029> A_IWL<21028> A_IWL<21027> A_IWL<21026> A_IWL<21025> A_IWL<21024> A_IWL<21023> A_IWL<21022> A_IWL<21021> A_IWL<21020> A_IWL<21019> A_IWL<21018> A_IWL<21017> A_IWL<21016> A_IWL<21015> A_IWL<21014> A_IWL<21013> A_IWL<21012> A_IWL<21011> A_IWL<21010> A_IWL<21009> A_IWL<21008> A_IWL<21007> A_IWL<21006> A_IWL<21005> A_IWL<21004> A_IWL<21003> A_IWL<21002> A_IWL<21001> A_IWL<21000> A_IWL<20999> A_IWL<20998> A_IWL<20997> A_IWL<20996> A_IWL<20995> A_IWL<20994> A_IWL<20993> A_IWL<20992> A_IWL<22015> A_IWL<22014> A_IWL<22013> A_IWL<22012> A_IWL<22011> A_IWL<22010> A_IWL<22009> A_IWL<22008> A_IWL<22007> A_IWL<22006> A_IWL<22005> A_IWL<22004> A_IWL<22003> A_IWL<22002> A_IWL<22001> A_IWL<22000> A_IWL<21999> A_IWL<21998> A_IWL<21997> A_IWL<21996> A_IWL<21995> A_IWL<21994> A_IWL<21993> A_IWL<21992> A_IWL<21991> A_IWL<21990> A_IWL<21989> A_IWL<21988> A_IWL<21987> A_IWL<21986> A_IWL<21985> A_IWL<21984> A_IWL<21983> A_IWL<21982> A_IWL<21981> A_IWL<21980> A_IWL<21979> A_IWL<21978> A_IWL<21977> A_IWL<21976> A_IWL<21975> A_IWL<21974> A_IWL<21973> A_IWL<21972> A_IWL<21971> A_IWL<21970> A_IWL<21969> A_IWL<21968> A_IWL<21967> A_IWL<21966> A_IWL<21965> A_IWL<21964> A_IWL<21963> A_IWL<21962> A_IWL<21961> A_IWL<21960> A_IWL<21959> A_IWL<21958> A_IWL<21957> A_IWL<21956> A_IWL<21955> A_IWL<21954> A_IWL<21953> A_IWL<21952> A_IWL<21951> A_IWL<21950> A_IWL<21949> A_IWL<21948> A_IWL<21947> A_IWL<21946> A_IWL<21945> A_IWL<21944> A_IWL<21943> A_IWL<21942> A_IWL<21941> A_IWL<21940> A_IWL<21939> A_IWL<21938> A_IWL<21937> A_IWL<21936> A_IWL<21935> A_IWL<21934> A_IWL<21933> A_IWL<21932> A_IWL<21931> A_IWL<21930> A_IWL<21929> A_IWL<21928> A_IWL<21927> A_IWL<21926> A_IWL<21925> A_IWL<21924> A_IWL<21923> A_IWL<21922> A_IWL<21921> A_IWL<21920> A_IWL<21919> A_IWL<21918> A_IWL<21917> A_IWL<21916> A_IWL<21915> A_IWL<21914> A_IWL<21913> A_IWL<21912> A_IWL<21911> A_IWL<21910> A_IWL<21909> A_IWL<21908> A_IWL<21907> A_IWL<21906> A_IWL<21905> A_IWL<21904> A_IWL<21903> A_IWL<21902> A_IWL<21901> A_IWL<21900> A_IWL<21899> A_IWL<21898> A_IWL<21897> A_IWL<21896> A_IWL<21895> A_IWL<21894> A_IWL<21893> A_IWL<21892> A_IWL<21891> A_IWL<21890> A_IWL<21889> A_IWL<21888> A_IWL<21887> A_IWL<21886> A_IWL<21885> A_IWL<21884> A_IWL<21883> A_IWL<21882> A_IWL<21881> A_IWL<21880> A_IWL<21879> A_IWL<21878> A_IWL<21877> A_IWL<21876> A_IWL<21875> A_IWL<21874> A_IWL<21873> A_IWL<21872> A_IWL<21871> A_IWL<21870> A_IWL<21869> A_IWL<21868> A_IWL<21867> A_IWL<21866> A_IWL<21865> A_IWL<21864> A_IWL<21863> A_IWL<21862> A_IWL<21861> A_IWL<21860> A_IWL<21859> A_IWL<21858> A_IWL<21857> A_IWL<21856> A_IWL<21855> A_IWL<21854> A_IWL<21853> A_IWL<21852> A_IWL<21851> A_IWL<21850> A_IWL<21849> A_IWL<21848> A_IWL<21847> A_IWL<21846> A_IWL<21845> A_IWL<21844> A_IWL<21843> A_IWL<21842> A_IWL<21841> A_IWL<21840> A_IWL<21839> A_IWL<21838> A_IWL<21837> A_IWL<21836> A_IWL<21835> A_IWL<21834> A_IWL<21833> A_IWL<21832> A_IWL<21831> A_IWL<21830> A_IWL<21829> A_IWL<21828> A_IWL<21827> A_IWL<21826> A_IWL<21825> A_IWL<21824> A_IWL<21823> A_IWL<21822> A_IWL<21821> A_IWL<21820> A_IWL<21819> A_IWL<21818> A_IWL<21817> A_IWL<21816> A_IWL<21815> A_IWL<21814> A_IWL<21813> A_IWL<21812> A_IWL<21811> A_IWL<21810> A_IWL<21809> A_IWL<21808> A_IWL<21807> A_IWL<21806> A_IWL<21805> A_IWL<21804> A_IWL<21803> A_IWL<21802> A_IWL<21801> A_IWL<21800> A_IWL<21799> A_IWL<21798> A_IWL<21797> A_IWL<21796> A_IWL<21795> A_IWL<21794> A_IWL<21793> A_IWL<21792> A_IWL<21791> A_IWL<21790> A_IWL<21789> A_IWL<21788> A_IWL<21787> A_IWL<21786> A_IWL<21785> A_IWL<21784> A_IWL<21783> A_IWL<21782> A_IWL<21781> A_IWL<21780> A_IWL<21779> A_IWL<21778> A_IWL<21777> A_IWL<21776> A_IWL<21775> A_IWL<21774> A_IWL<21773> A_IWL<21772> A_IWL<21771> A_IWL<21770> A_IWL<21769> A_IWL<21768> A_IWL<21767> A_IWL<21766> A_IWL<21765> A_IWL<21764> A_IWL<21763> A_IWL<21762> A_IWL<21761> A_IWL<21760> A_IWL<21759> A_IWL<21758> A_IWL<21757> A_IWL<21756> A_IWL<21755> A_IWL<21754> A_IWL<21753> A_IWL<21752> A_IWL<21751> A_IWL<21750> A_IWL<21749> A_IWL<21748> A_IWL<21747> A_IWL<21746> A_IWL<21745> A_IWL<21744> A_IWL<21743> A_IWL<21742> A_IWL<21741> A_IWL<21740> A_IWL<21739> A_IWL<21738> A_IWL<21737> A_IWL<21736> A_IWL<21735> A_IWL<21734> A_IWL<21733> A_IWL<21732> A_IWL<21731> A_IWL<21730> A_IWL<21729> A_IWL<21728> A_IWL<21727> A_IWL<21726> A_IWL<21725> A_IWL<21724> A_IWL<21723> A_IWL<21722> A_IWL<21721> A_IWL<21720> A_IWL<21719> A_IWL<21718> A_IWL<21717> A_IWL<21716> A_IWL<21715> A_IWL<21714> A_IWL<21713> A_IWL<21712> A_IWL<21711> A_IWL<21710> A_IWL<21709> A_IWL<21708> A_IWL<21707> A_IWL<21706> A_IWL<21705> A_IWL<21704> A_IWL<21703> A_IWL<21702> A_IWL<21701> A_IWL<21700> A_IWL<21699> A_IWL<21698> A_IWL<21697> A_IWL<21696> A_IWL<21695> A_IWL<21694> A_IWL<21693> A_IWL<21692> A_IWL<21691> A_IWL<21690> A_IWL<21689> A_IWL<21688> A_IWL<21687> A_IWL<21686> A_IWL<21685> A_IWL<21684> A_IWL<21683> A_IWL<21682> A_IWL<21681> A_IWL<21680> A_IWL<21679> A_IWL<21678> A_IWL<21677> A_IWL<21676> A_IWL<21675> A_IWL<21674> A_IWL<21673> A_IWL<21672> A_IWL<21671> A_IWL<21670> A_IWL<21669> A_IWL<21668> A_IWL<21667> A_IWL<21666> A_IWL<21665> A_IWL<21664> A_IWL<21663> A_IWL<21662> A_IWL<21661> A_IWL<21660> A_IWL<21659> A_IWL<21658> A_IWL<21657> A_IWL<21656> A_IWL<21655> A_IWL<21654> A_IWL<21653> A_IWL<21652> A_IWL<21651> A_IWL<21650> A_IWL<21649> A_IWL<21648> A_IWL<21647> A_IWL<21646> A_IWL<21645> A_IWL<21644> A_IWL<21643> A_IWL<21642> A_IWL<21641> A_IWL<21640> A_IWL<21639> A_IWL<21638> A_IWL<21637> A_IWL<21636> A_IWL<21635> A_IWL<21634> A_IWL<21633> A_IWL<21632> A_IWL<21631> A_IWL<21630> A_IWL<21629> A_IWL<21628> A_IWL<21627> A_IWL<21626> A_IWL<21625> A_IWL<21624> A_IWL<21623> A_IWL<21622> A_IWL<21621> A_IWL<21620> A_IWL<21619> A_IWL<21618> A_IWL<21617> A_IWL<21616> A_IWL<21615> A_IWL<21614> A_IWL<21613> A_IWL<21612> A_IWL<21611> A_IWL<21610> A_IWL<21609> A_IWL<21608> A_IWL<21607> A_IWL<21606> A_IWL<21605> A_IWL<21604> A_IWL<21603> A_IWL<21602> A_IWL<21601> A_IWL<21600> A_IWL<21599> A_IWL<21598> A_IWL<21597> A_IWL<21596> A_IWL<21595> A_IWL<21594> A_IWL<21593> A_IWL<21592> A_IWL<21591> A_IWL<21590> A_IWL<21589> A_IWL<21588> A_IWL<21587> A_IWL<21586> A_IWL<21585> A_IWL<21584> A_IWL<21583> A_IWL<21582> A_IWL<21581> A_IWL<21580> A_IWL<21579> A_IWL<21578> A_IWL<21577> A_IWL<21576> A_IWL<21575> A_IWL<21574> A_IWL<21573> A_IWL<21572> A_IWL<21571> A_IWL<21570> A_IWL<21569> A_IWL<21568> A_IWL<21567> A_IWL<21566> A_IWL<21565> A_IWL<21564> A_IWL<21563> A_IWL<21562> A_IWL<21561> A_IWL<21560> A_IWL<21559> A_IWL<21558> A_IWL<21557> A_IWL<21556> A_IWL<21555> A_IWL<21554> A_IWL<21553> A_IWL<21552> A_IWL<21551> A_IWL<21550> A_IWL<21549> A_IWL<21548> A_IWL<21547> A_IWL<21546> A_IWL<21545> A_IWL<21544> A_IWL<21543> A_IWL<21542> A_IWL<21541> A_IWL<21540> A_IWL<21539> A_IWL<21538> A_IWL<21537> A_IWL<21536> A_IWL<21535> A_IWL<21534> A_IWL<21533> A_IWL<21532> A_IWL<21531> A_IWL<21530> A_IWL<21529> A_IWL<21528> A_IWL<21527> A_IWL<21526> A_IWL<21525> A_IWL<21524> A_IWL<21523> A_IWL<21522> A_IWL<21521> A_IWL<21520> A_IWL<21519> A_IWL<21518> A_IWL<21517> A_IWL<21516> A_IWL<21515> A_IWL<21514> A_IWL<21513> A_IWL<21512> A_IWL<21511> A_IWL<21510> A_IWL<21509> A_IWL<21508> A_IWL<21507> A_IWL<21506> A_IWL<21505> A_IWL<21504> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<41> A_BLC<83> A_BLC<82> A_BLC_TOP<83> A_BLC_TOP<82> A_BLT<83> A_BLT<82> A_BLT_TOP<83> A_BLT_TOP<82> A_IWL<20991> A_IWL<20990> A_IWL<20989> A_IWL<20988> A_IWL<20987> A_IWL<20986> A_IWL<20985> A_IWL<20984> A_IWL<20983> A_IWL<20982> A_IWL<20981> A_IWL<20980> A_IWL<20979> A_IWL<20978> A_IWL<20977> A_IWL<20976> A_IWL<20975> A_IWL<20974> A_IWL<20973> A_IWL<20972> A_IWL<20971> A_IWL<20970> A_IWL<20969> A_IWL<20968> A_IWL<20967> A_IWL<20966> A_IWL<20965> A_IWL<20964> A_IWL<20963> A_IWL<20962> A_IWL<20961> A_IWL<20960> A_IWL<20959> A_IWL<20958> A_IWL<20957> A_IWL<20956> A_IWL<20955> A_IWL<20954> A_IWL<20953> A_IWL<20952> A_IWL<20951> A_IWL<20950> A_IWL<20949> A_IWL<20948> A_IWL<20947> A_IWL<20946> A_IWL<20945> A_IWL<20944> A_IWL<20943> A_IWL<20942> A_IWL<20941> A_IWL<20940> A_IWL<20939> A_IWL<20938> A_IWL<20937> A_IWL<20936> A_IWL<20935> A_IWL<20934> A_IWL<20933> A_IWL<20932> A_IWL<20931> A_IWL<20930> A_IWL<20929> A_IWL<20928> A_IWL<20927> A_IWL<20926> A_IWL<20925> A_IWL<20924> A_IWL<20923> A_IWL<20922> A_IWL<20921> A_IWL<20920> A_IWL<20919> A_IWL<20918> A_IWL<20917> A_IWL<20916> A_IWL<20915> A_IWL<20914> A_IWL<20913> A_IWL<20912> A_IWL<20911> A_IWL<20910> A_IWL<20909> A_IWL<20908> A_IWL<20907> A_IWL<20906> A_IWL<20905> A_IWL<20904> A_IWL<20903> A_IWL<20902> A_IWL<20901> A_IWL<20900> A_IWL<20899> A_IWL<20898> A_IWL<20897> A_IWL<20896> A_IWL<20895> A_IWL<20894> A_IWL<20893> A_IWL<20892> A_IWL<20891> A_IWL<20890> A_IWL<20889> A_IWL<20888> A_IWL<20887> A_IWL<20886> A_IWL<20885> A_IWL<20884> A_IWL<20883> A_IWL<20882> A_IWL<20881> A_IWL<20880> A_IWL<20879> A_IWL<20878> A_IWL<20877> A_IWL<20876> A_IWL<20875> A_IWL<20874> A_IWL<20873> A_IWL<20872> A_IWL<20871> A_IWL<20870> A_IWL<20869> A_IWL<20868> A_IWL<20867> A_IWL<20866> A_IWL<20865> A_IWL<20864> A_IWL<20863> A_IWL<20862> A_IWL<20861> A_IWL<20860> A_IWL<20859> A_IWL<20858> A_IWL<20857> A_IWL<20856> A_IWL<20855> A_IWL<20854> A_IWL<20853> A_IWL<20852> A_IWL<20851> A_IWL<20850> A_IWL<20849> A_IWL<20848> A_IWL<20847> A_IWL<20846> A_IWL<20845> A_IWL<20844> A_IWL<20843> A_IWL<20842> A_IWL<20841> A_IWL<20840> A_IWL<20839> A_IWL<20838> A_IWL<20837> A_IWL<20836> A_IWL<20835> A_IWL<20834> A_IWL<20833> A_IWL<20832> A_IWL<20831> A_IWL<20830> A_IWL<20829> A_IWL<20828> A_IWL<20827> A_IWL<20826> A_IWL<20825> A_IWL<20824> A_IWL<20823> A_IWL<20822> A_IWL<20821> A_IWL<20820> A_IWL<20819> A_IWL<20818> A_IWL<20817> A_IWL<20816> A_IWL<20815> A_IWL<20814> A_IWL<20813> A_IWL<20812> A_IWL<20811> A_IWL<20810> A_IWL<20809> A_IWL<20808> A_IWL<20807> A_IWL<20806> A_IWL<20805> A_IWL<20804> A_IWL<20803> A_IWL<20802> A_IWL<20801> A_IWL<20800> A_IWL<20799> A_IWL<20798> A_IWL<20797> A_IWL<20796> A_IWL<20795> A_IWL<20794> A_IWL<20793> A_IWL<20792> A_IWL<20791> A_IWL<20790> A_IWL<20789> A_IWL<20788> A_IWL<20787> A_IWL<20786> A_IWL<20785> A_IWL<20784> A_IWL<20783> A_IWL<20782> A_IWL<20781> A_IWL<20780> A_IWL<20779> A_IWL<20778> A_IWL<20777> A_IWL<20776> A_IWL<20775> A_IWL<20774> A_IWL<20773> A_IWL<20772> A_IWL<20771> A_IWL<20770> A_IWL<20769> A_IWL<20768> A_IWL<20767> A_IWL<20766> A_IWL<20765> A_IWL<20764> A_IWL<20763> A_IWL<20762> A_IWL<20761> A_IWL<20760> A_IWL<20759> A_IWL<20758> A_IWL<20757> A_IWL<20756> A_IWL<20755> A_IWL<20754> A_IWL<20753> A_IWL<20752> A_IWL<20751> A_IWL<20750> A_IWL<20749> A_IWL<20748> A_IWL<20747> A_IWL<20746> A_IWL<20745> A_IWL<20744> A_IWL<20743> A_IWL<20742> A_IWL<20741> A_IWL<20740> A_IWL<20739> A_IWL<20738> A_IWL<20737> A_IWL<20736> A_IWL<20735> A_IWL<20734> A_IWL<20733> A_IWL<20732> A_IWL<20731> A_IWL<20730> A_IWL<20729> A_IWL<20728> A_IWL<20727> A_IWL<20726> A_IWL<20725> A_IWL<20724> A_IWL<20723> A_IWL<20722> A_IWL<20721> A_IWL<20720> A_IWL<20719> A_IWL<20718> A_IWL<20717> A_IWL<20716> A_IWL<20715> A_IWL<20714> A_IWL<20713> A_IWL<20712> A_IWL<20711> A_IWL<20710> A_IWL<20709> A_IWL<20708> A_IWL<20707> A_IWL<20706> A_IWL<20705> A_IWL<20704> A_IWL<20703> A_IWL<20702> A_IWL<20701> A_IWL<20700> A_IWL<20699> A_IWL<20698> A_IWL<20697> A_IWL<20696> A_IWL<20695> A_IWL<20694> A_IWL<20693> A_IWL<20692> A_IWL<20691> A_IWL<20690> A_IWL<20689> A_IWL<20688> A_IWL<20687> A_IWL<20686> A_IWL<20685> A_IWL<20684> A_IWL<20683> A_IWL<20682> A_IWL<20681> A_IWL<20680> A_IWL<20679> A_IWL<20678> A_IWL<20677> A_IWL<20676> A_IWL<20675> A_IWL<20674> A_IWL<20673> A_IWL<20672> A_IWL<20671> A_IWL<20670> A_IWL<20669> A_IWL<20668> A_IWL<20667> A_IWL<20666> A_IWL<20665> A_IWL<20664> A_IWL<20663> A_IWL<20662> A_IWL<20661> A_IWL<20660> A_IWL<20659> A_IWL<20658> A_IWL<20657> A_IWL<20656> A_IWL<20655> A_IWL<20654> A_IWL<20653> A_IWL<20652> A_IWL<20651> A_IWL<20650> A_IWL<20649> A_IWL<20648> A_IWL<20647> A_IWL<20646> A_IWL<20645> A_IWL<20644> A_IWL<20643> A_IWL<20642> A_IWL<20641> A_IWL<20640> A_IWL<20639> A_IWL<20638> A_IWL<20637> A_IWL<20636> A_IWL<20635> A_IWL<20634> A_IWL<20633> A_IWL<20632> A_IWL<20631> A_IWL<20630> A_IWL<20629> A_IWL<20628> A_IWL<20627> A_IWL<20626> A_IWL<20625> A_IWL<20624> A_IWL<20623> A_IWL<20622> A_IWL<20621> A_IWL<20620> A_IWL<20619> A_IWL<20618> A_IWL<20617> A_IWL<20616> A_IWL<20615> A_IWL<20614> A_IWL<20613> A_IWL<20612> A_IWL<20611> A_IWL<20610> A_IWL<20609> A_IWL<20608> A_IWL<20607> A_IWL<20606> A_IWL<20605> A_IWL<20604> A_IWL<20603> A_IWL<20602> A_IWL<20601> A_IWL<20600> A_IWL<20599> A_IWL<20598> A_IWL<20597> A_IWL<20596> A_IWL<20595> A_IWL<20594> A_IWL<20593> A_IWL<20592> A_IWL<20591> A_IWL<20590> A_IWL<20589> A_IWL<20588> A_IWL<20587> A_IWL<20586> A_IWL<20585> A_IWL<20584> A_IWL<20583> A_IWL<20582> A_IWL<20581> A_IWL<20580> A_IWL<20579> A_IWL<20578> A_IWL<20577> A_IWL<20576> A_IWL<20575> A_IWL<20574> A_IWL<20573> A_IWL<20572> A_IWL<20571> A_IWL<20570> A_IWL<20569> A_IWL<20568> A_IWL<20567> A_IWL<20566> A_IWL<20565> A_IWL<20564> A_IWL<20563> A_IWL<20562> A_IWL<20561> A_IWL<20560> A_IWL<20559> A_IWL<20558> A_IWL<20557> A_IWL<20556> A_IWL<20555> A_IWL<20554> A_IWL<20553> A_IWL<20552> A_IWL<20551> A_IWL<20550> A_IWL<20549> A_IWL<20548> A_IWL<20547> A_IWL<20546> A_IWL<20545> A_IWL<20544> A_IWL<20543> A_IWL<20542> A_IWL<20541> A_IWL<20540> A_IWL<20539> A_IWL<20538> A_IWL<20537> A_IWL<20536> A_IWL<20535> A_IWL<20534> A_IWL<20533> A_IWL<20532> A_IWL<20531> A_IWL<20530> A_IWL<20529> A_IWL<20528> A_IWL<20527> A_IWL<20526> A_IWL<20525> A_IWL<20524> A_IWL<20523> A_IWL<20522> A_IWL<20521> A_IWL<20520> A_IWL<20519> A_IWL<20518> A_IWL<20517> A_IWL<20516> A_IWL<20515> A_IWL<20514> A_IWL<20513> A_IWL<20512> A_IWL<20511> A_IWL<20510> A_IWL<20509> A_IWL<20508> A_IWL<20507> A_IWL<20506> A_IWL<20505> A_IWL<20504> A_IWL<20503> A_IWL<20502> A_IWL<20501> A_IWL<20500> A_IWL<20499> A_IWL<20498> A_IWL<20497> A_IWL<20496> A_IWL<20495> A_IWL<20494> A_IWL<20493> A_IWL<20492> A_IWL<20491> A_IWL<20490> A_IWL<20489> A_IWL<20488> A_IWL<20487> A_IWL<20486> A_IWL<20485> A_IWL<20484> A_IWL<20483> A_IWL<20482> A_IWL<20481> A_IWL<20480> A_IWL<21503> A_IWL<21502> A_IWL<21501> A_IWL<21500> A_IWL<21499> A_IWL<21498> A_IWL<21497> A_IWL<21496> A_IWL<21495> A_IWL<21494> A_IWL<21493> A_IWL<21492> A_IWL<21491> A_IWL<21490> A_IWL<21489> A_IWL<21488> A_IWL<21487> A_IWL<21486> A_IWL<21485> A_IWL<21484> A_IWL<21483> A_IWL<21482> A_IWL<21481> A_IWL<21480> A_IWL<21479> A_IWL<21478> A_IWL<21477> A_IWL<21476> A_IWL<21475> A_IWL<21474> A_IWL<21473> A_IWL<21472> A_IWL<21471> A_IWL<21470> A_IWL<21469> A_IWL<21468> A_IWL<21467> A_IWL<21466> A_IWL<21465> A_IWL<21464> A_IWL<21463> A_IWL<21462> A_IWL<21461> A_IWL<21460> A_IWL<21459> A_IWL<21458> A_IWL<21457> A_IWL<21456> A_IWL<21455> A_IWL<21454> A_IWL<21453> A_IWL<21452> A_IWL<21451> A_IWL<21450> A_IWL<21449> A_IWL<21448> A_IWL<21447> A_IWL<21446> A_IWL<21445> A_IWL<21444> A_IWL<21443> A_IWL<21442> A_IWL<21441> A_IWL<21440> A_IWL<21439> A_IWL<21438> A_IWL<21437> A_IWL<21436> A_IWL<21435> A_IWL<21434> A_IWL<21433> A_IWL<21432> A_IWL<21431> A_IWL<21430> A_IWL<21429> A_IWL<21428> A_IWL<21427> A_IWL<21426> A_IWL<21425> A_IWL<21424> A_IWL<21423> A_IWL<21422> A_IWL<21421> A_IWL<21420> A_IWL<21419> A_IWL<21418> A_IWL<21417> A_IWL<21416> A_IWL<21415> A_IWL<21414> A_IWL<21413> A_IWL<21412> A_IWL<21411> A_IWL<21410> A_IWL<21409> A_IWL<21408> A_IWL<21407> A_IWL<21406> A_IWL<21405> A_IWL<21404> A_IWL<21403> A_IWL<21402> A_IWL<21401> A_IWL<21400> A_IWL<21399> A_IWL<21398> A_IWL<21397> A_IWL<21396> A_IWL<21395> A_IWL<21394> A_IWL<21393> A_IWL<21392> A_IWL<21391> A_IWL<21390> A_IWL<21389> A_IWL<21388> A_IWL<21387> A_IWL<21386> A_IWL<21385> A_IWL<21384> A_IWL<21383> A_IWL<21382> A_IWL<21381> A_IWL<21380> A_IWL<21379> A_IWL<21378> A_IWL<21377> A_IWL<21376> A_IWL<21375> A_IWL<21374> A_IWL<21373> A_IWL<21372> A_IWL<21371> A_IWL<21370> A_IWL<21369> A_IWL<21368> A_IWL<21367> A_IWL<21366> A_IWL<21365> A_IWL<21364> A_IWL<21363> A_IWL<21362> A_IWL<21361> A_IWL<21360> A_IWL<21359> A_IWL<21358> A_IWL<21357> A_IWL<21356> A_IWL<21355> A_IWL<21354> A_IWL<21353> A_IWL<21352> A_IWL<21351> A_IWL<21350> A_IWL<21349> A_IWL<21348> A_IWL<21347> A_IWL<21346> A_IWL<21345> A_IWL<21344> A_IWL<21343> A_IWL<21342> A_IWL<21341> A_IWL<21340> A_IWL<21339> A_IWL<21338> A_IWL<21337> A_IWL<21336> A_IWL<21335> A_IWL<21334> A_IWL<21333> A_IWL<21332> A_IWL<21331> A_IWL<21330> A_IWL<21329> A_IWL<21328> A_IWL<21327> A_IWL<21326> A_IWL<21325> A_IWL<21324> A_IWL<21323> A_IWL<21322> A_IWL<21321> A_IWL<21320> A_IWL<21319> A_IWL<21318> A_IWL<21317> A_IWL<21316> A_IWL<21315> A_IWL<21314> A_IWL<21313> A_IWL<21312> A_IWL<21311> A_IWL<21310> A_IWL<21309> A_IWL<21308> A_IWL<21307> A_IWL<21306> A_IWL<21305> A_IWL<21304> A_IWL<21303> A_IWL<21302> A_IWL<21301> A_IWL<21300> A_IWL<21299> A_IWL<21298> A_IWL<21297> A_IWL<21296> A_IWL<21295> A_IWL<21294> A_IWL<21293> A_IWL<21292> A_IWL<21291> A_IWL<21290> A_IWL<21289> A_IWL<21288> A_IWL<21287> A_IWL<21286> A_IWL<21285> A_IWL<21284> A_IWL<21283> A_IWL<21282> A_IWL<21281> A_IWL<21280> A_IWL<21279> A_IWL<21278> A_IWL<21277> A_IWL<21276> A_IWL<21275> A_IWL<21274> A_IWL<21273> A_IWL<21272> A_IWL<21271> A_IWL<21270> A_IWL<21269> A_IWL<21268> A_IWL<21267> A_IWL<21266> A_IWL<21265> A_IWL<21264> A_IWL<21263> A_IWL<21262> A_IWL<21261> A_IWL<21260> A_IWL<21259> A_IWL<21258> A_IWL<21257> A_IWL<21256> A_IWL<21255> A_IWL<21254> A_IWL<21253> A_IWL<21252> A_IWL<21251> A_IWL<21250> A_IWL<21249> A_IWL<21248> A_IWL<21247> A_IWL<21246> A_IWL<21245> A_IWL<21244> A_IWL<21243> A_IWL<21242> A_IWL<21241> A_IWL<21240> A_IWL<21239> A_IWL<21238> A_IWL<21237> A_IWL<21236> A_IWL<21235> A_IWL<21234> A_IWL<21233> A_IWL<21232> A_IWL<21231> A_IWL<21230> A_IWL<21229> A_IWL<21228> A_IWL<21227> A_IWL<21226> A_IWL<21225> A_IWL<21224> A_IWL<21223> A_IWL<21222> A_IWL<21221> A_IWL<21220> A_IWL<21219> A_IWL<21218> A_IWL<21217> A_IWL<21216> A_IWL<21215> A_IWL<21214> A_IWL<21213> A_IWL<21212> A_IWL<21211> A_IWL<21210> A_IWL<21209> A_IWL<21208> A_IWL<21207> A_IWL<21206> A_IWL<21205> A_IWL<21204> A_IWL<21203> A_IWL<21202> A_IWL<21201> A_IWL<21200> A_IWL<21199> A_IWL<21198> A_IWL<21197> A_IWL<21196> A_IWL<21195> A_IWL<21194> A_IWL<21193> A_IWL<21192> A_IWL<21191> A_IWL<21190> A_IWL<21189> A_IWL<21188> A_IWL<21187> A_IWL<21186> A_IWL<21185> A_IWL<21184> A_IWL<21183> A_IWL<21182> A_IWL<21181> A_IWL<21180> A_IWL<21179> A_IWL<21178> A_IWL<21177> A_IWL<21176> A_IWL<21175> A_IWL<21174> A_IWL<21173> A_IWL<21172> A_IWL<21171> A_IWL<21170> A_IWL<21169> A_IWL<21168> A_IWL<21167> A_IWL<21166> A_IWL<21165> A_IWL<21164> A_IWL<21163> A_IWL<21162> A_IWL<21161> A_IWL<21160> A_IWL<21159> A_IWL<21158> A_IWL<21157> A_IWL<21156> A_IWL<21155> A_IWL<21154> A_IWL<21153> A_IWL<21152> A_IWL<21151> A_IWL<21150> A_IWL<21149> A_IWL<21148> A_IWL<21147> A_IWL<21146> A_IWL<21145> A_IWL<21144> A_IWL<21143> A_IWL<21142> A_IWL<21141> A_IWL<21140> A_IWL<21139> A_IWL<21138> A_IWL<21137> A_IWL<21136> A_IWL<21135> A_IWL<21134> A_IWL<21133> A_IWL<21132> A_IWL<21131> A_IWL<21130> A_IWL<21129> A_IWL<21128> A_IWL<21127> A_IWL<21126> A_IWL<21125> A_IWL<21124> A_IWL<21123> A_IWL<21122> A_IWL<21121> A_IWL<21120> A_IWL<21119> A_IWL<21118> A_IWL<21117> A_IWL<21116> A_IWL<21115> A_IWL<21114> A_IWL<21113> A_IWL<21112> A_IWL<21111> A_IWL<21110> A_IWL<21109> A_IWL<21108> A_IWL<21107> A_IWL<21106> A_IWL<21105> A_IWL<21104> A_IWL<21103> A_IWL<21102> A_IWL<21101> A_IWL<21100> A_IWL<21099> A_IWL<21098> A_IWL<21097> A_IWL<21096> A_IWL<21095> A_IWL<21094> A_IWL<21093> A_IWL<21092> A_IWL<21091> A_IWL<21090> A_IWL<21089> A_IWL<21088> A_IWL<21087> A_IWL<21086> A_IWL<21085> A_IWL<21084> A_IWL<21083> A_IWL<21082> A_IWL<21081> A_IWL<21080> A_IWL<21079> A_IWL<21078> A_IWL<21077> A_IWL<21076> A_IWL<21075> A_IWL<21074> A_IWL<21073> A_IWL<21072> A_IWL<21071> A_IWL<21070> A_IWL<21069> A_IWL<21068> A_IWL<21067> A_IWL<21066> A_IWL<21065> A_IWL<21064> A_IWL<21063> A_IWL<21062> A_IWL<21061> A_IWL<21060> A_IWL<21059> A_IWL<21058> A_IWL<21057> A_IWL<21056> A_IWL<21055> A_IWL<21054> A_IWL<21053> A_IWL<21052> A_IWL<21051> A_IWL<21050> A_IWL<21049> A_IWL<21048> A_IWL<21047> A_IWL<21046> A_IWL<21045> A_IWL<21044> A_IWL<21043> A_IWL<21042> A_IWL<21041> A_IWL<21040> A_IWL<21039> A_IWL<21038> A_IWL<21037> A_IWL<21036> A_IWL<21035> A_IWL<21034> A_IWL<21033> A_IWL<21032> A_IWL<21031> A_IWL<21030> A_IWL<21029> A_IWL<21028> A_IWL<21027> A_IWL<21026> A_IWL<21025> A_IWL<21024> A_IWL<21023> A_IWL<21022> A_IWL<21021> A_IWL<21020> A_IWL<21019> A_IWL<21018> A_IWL<21017> A_IWL<21016> A_IWL<21015> A_IWL<21014> A_IWL<21013> A_IWL<21012> A_IWL<21011> A_IWL<21010> A_IWL<21009> A_IWL<21008> A_IWL<21007> A_IWL<21006> A_IWL<21005> A_IWL<21004> A_IWL<21003> A_IWL<21002> A_IWL<21001> A_IWL<21000> A_IWL<20999> A_IWL<20998> A_IWL<20997> A_IWL<20996> A_IWL<20995> A_IWL<20994> A_IWL<20993> A_IWL<20992> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<40> A_BLC<81> A_BLC<80> A_BLC_TOP<81> A_BLC_TOP<80> A_BLT<81> A_BLT<80> A_BLT_TOP<81> A_BLT_TOP<80> A_IWL<20479> A_IWL<20478> A_IWL<20477> A_IWL<20476> A_IWL<20475> A_IWL<20474> A_IWL<20473> A_IWL<20472> A_IWL<20471> A_IWL<20470> A_IWL<20469> A_IWL<20468> A_IWL<20467> A_IWL<20466> A_IWL<20465> A_IWL<20464> A_IWL<20463> A_IWL<20462> A_IWL<20461> A_IWL<20460> A_IWL<20459> A_IWL<20458> A_IWL<20457> A_IWL<20456> A_IWL<20455> A_IWL<20454> A_IWL<20453> A_IWL<20452> A_IWL<20451> A_IWL<20450> A_IWL<20449> A_IWL<20448> A_IWL<20447> A_IWL<20446> A_IWL<20445> A_IWL<20444> A_IWL<20443> A_IWL<20442> A_IWL<20441> A_IWL<20440> A_IWL<20439> A_IWL<20438> A_IWL<20437> A_IWL<20436> A_IWL<20435> A_IWL<20434> A_IWL<20433> A_IWL<20432> A_IWL<20431> A_IWL<20430> A_IWL<20429> A_IWL<20428> A_IWL<20427> A_IWL<20426> A_IWL<20425> A_IWL<20424> A_IWL<20423> A_IWL<20422> A_IWL<20421> A_IWL<20420> A_IWL<20419> A_IWL<20418> A_IWL<20417> A_IWL<20416> A_IWL<20415> A_IWL<20414> A_IWL<20413> A_IWL<20412> A_IWL<20411> A_IWL<20410> A_IWL<20409> A_IWL<20408> A_IWL<20407> A_IWL<20406> A_IWL<20405> A_IWL<20404> A_IWL<20403> A_IWL<20402> A_IWL<20401> A_IWL<20400> A_IWL<20399> A_IWL<20398> A_IWL<20397> A_IWL<20396> A_IWL<20395> A_IWL<20394> A_IWL<20393> A_IWL<20392> A_IWL<20391> A_IWL<20390> A_IWL<20389> A_IWL<20388> A_IWL<20387> A_IWL<20386> A_IWL<20385> A_IWL<20384> A_IWL<20383> A_IWL<20382> A_IWL<20381> A_IWL<20380> A_IWL<20379> A_IWL<20378> A_IWL<20377> A_IWL<20376> A_IWL<20375> A_IWL<20374> A_IWL<20373> A_IWL<20372> A_IWL<20371> A_IWL<20370> A_IWL<20369> A_IWL<20368> A_IWL<20367> A_IWL<20366> A_IWL<20365> A_IWL<20364> A_IWL<20363> A_IWL<20362> A_IWL<20361> A_IWL<20360> A_IWL<20359> A_IWL<20358> A_IWL<20357> A_IWL<20356> A_IWL<20355> A_IWL<20354> A_IWL<20353> A_IWL<20352> A_IWL<20351> A_IWL<20350> A_IWL<20349> A_IWL<20348> A_IWL<20347> A_IWL<20346> A_IWL<20345> A_IWL<20344> A_IWL<20343> A_IWL<20342> A_IWL<20341> A_IWL<20340> A_IWL<20339> A_IWL<20338> A_IWL<20337> A_IWL<20336> A_IWL<20335> A_IWL<20334> A_IWL<20333> A_IWL<20332> A_IWL<20331> A_IWL<20330> A_IWL<20329> A_IWL<20328> A_IWL<20327> A_IWL<20326> A_IWL<20325> A_IWL<20324> A_IWL<20323> A_IWL<20322> A_IWL<20321> A_IWL<20320> A_IWL<20319> A_IWL<20318> A_IWL<20317> A_IWL<20316> A_IWL<20315> A_IWL<20314> A_IWL<20313> A_IWL<20312> A_IWL<20311> A_IWL<20310> A_IWL<20309> A_IWL<20308> A_IWL<20307> A_IWL<20306> A_IWL<20305> A_IWL<20304> A_IWL<20303> A_IWL<20302> A_IWL<20301> A_IWL<20300> A_IWL<20299> A_IWL<20298> A_IWL<20297> A_IWL<20296> A_IWL<20295> A_IWL<20294> A_IWL<20293> A_IWL<20292> A_IWL<20291> A_IWL<20290> A_IWL<20289> A_IWL<20288> A_IWL<20287> A_IWL<20286> A_IWL<20285> A_IWL<20284> A_IWL<20283> A_IWL<20282> A_IWL<20281> A_IWL<20280> A_IWL<20279> A_IWL<20278> A_IWL<20277> A_IWL<20276> A_IWL<20275> A_IWL<20274> A_IWL<20273> A_IWL<20272> A_IWL<20271> A_IWL<20270> A_IWL<20269> A_IWL<20268> A_IWL<20267> A_IWL<20266> A_IWL<20265> A_IWL<20264> A_IWL<20263> A_IWL<20262> A_IWL<20261> A_IWL<20260> A_IWL<20259> A_IWL<20258> A_IWL<20257> A_IWL<20256> A_IWL<20255> A_IWL<20254> A_IWL<20253> A_IWL<20252> A_IWL<20251> A_IWL<20250> A_IWL<20249> A_IWL<20248> A_IWL<20247> A_IWL<20246> A_IWL<20245> A_IWL<20244> A_IWL<20243> A_IWL<20242> A_IWL<20241> A_IWL<20240> A_IWL<20239> A_IWL<20238> A_IWL<20237> A_IWL<20236> A_IWL<20235> A_IWL<20234> A_IWL<20233> A_IWL<20232> A_IWL<20231> A_IWL<20230> A_IWL<20229> A_IWL<20228> A_IWL<20227> A_IWL<20226> A_IWL<20225> A_IWL<20224> A_IWL<20223> A_IWL<20222> A_IWL<20221> A_IWL<20220> A_IWL<20219> A_IWL<20218> A_IWL<20217> A_IWL<20216> A_IWL<20215> A_IWL<20214> A_IWL<20213> A_IWL<20212> A_IWL<20211> A_IWL<20210> A_IWL<20209> A_IWL<20208> A_IWL<20207> A_IWL<20206> A_IWL<20205> A_IWL<20204> A_IWL<20203> A_IWL<20202> A_IWL<20201> A_IWL<20200> A_IWL<20199> A_IWL<20198> A_IWL<20197> A_IWL<20196> A_IWL<20195> A_IWL<20194> A_IWL<20193> A_IWL<20192> A_IWL<20191> A_IWL<20190> A_IWL<20189> A_IWL<20188> A_IWL<20187> A_IWL<20186> A_IWL<20185> A_IWL<20184> A_IWL<20183> A_IWL<20182> A_IWL<20181> A_IWL<20180> A_IWL<20179> A_IWL<20178> A_IWL<20177> A_IWL<20176> A_IWL<20175> A_IWL<20174> A_IWL<20173> A_IWL<20172> A_IWL<20171> A_IWL<20170> A_IWL<20169> A_IWL<20168> A_IWL<20167> A_IWL<20166> A_IWL<20165> A_IWL<20164> A_IWL<20163> A_IWL<20162> A_IWL<20161> A_IWL<20160> A_IWL<20159> A_IWL<20158> A_IWL<20157> A_IWL<20156> A_IWL<20155> A_IWL<20154> A_IWL<20153> A_IWL<20152> A_IWL<20151> A_IWL<20150> A_IWL<20149> A_IWL<20148> A_IWL<20147> A_IWL<20146> A_IWL<20145> A_IWL<20144> A_IWL<20143> A_IWL<20142> A_IWL<20141> A_IWL<20140> A_IWL<20139> A_IWL<20138> A_IWL<20137> A_IWL<20136> A_IWL<20135> A_IWL<20134> A_IWL<20133> A_IWL<20132> A_IWL<20131> A_IWL<20130> A_IWL<20129> A_IWL<20128> A_IWL<20127> A_IWL<20126> A_IWL<20125> A_IWL<20124> A_IWL<20123> A_IWL<20122> A_IWL<20121> A_IWL<20120> A_IWL<20119> A_IWL<20118> A_IWL<20117> A_IWL<20116> A_IWL<20115> A_IWL<20114> A_IWL<20113> A_IWL<20112> A_IWL<20111> A_IWL<20110> A_IWL<20109> A_IWL<20108> A_IWL<20107> A_IWL<20106> A_IWL<20105> A_IWL<20104> A_IWL<20103> A_IWL<20102> A_IWL<20101> A_IWL<20100> A_IWL<20099> A_IWL<20098> A_IWL<20097> A_IWL<20096> A_IWL<20095> A_IWL<20094> A_IWL<20093> A_IWL<20092> A_IWL<20091> A_IWL<20090> A_IWL<20089> A_IWL<20088> A_IWL<20087> A_IWL<20086> A_IWL<20085> A_IWL<20084> A_IWL<20083> A_IWL<20082> A_IWL<20081> A_IWL<20080> A_IWL<20079> A_IWL<20078> A_IWL<20077> A_IWL<20076> A_IWL<20075> A_IWL<20074> A_IWL<20073> A_IWL<20072> A_IWL<20071> A_IWL<20070> A_IWL<20069> A_IWL<20068> A_IWL<20067> A_IWL<20066> A_IWL<20065> A_IWL<20064> A_IWL<20063> A_IWL<20062> A_IWL<20061> A_IWL<20060> A_IWL<20059> A_IWL<20058> A_IWL<20057> A_IWL<20056> A_IWL<20055> A_IWL<20054> A_IWL<20053> A_IWL<20052> A_IWL<20051> A_IWL<20050> A_IWL<20049> A_IWL<20048> A_IWL<20047> A_IWL<20046> A_IWL<20045> A_IWL<20044> A_IWL<20043> A_IWL<20042> A_IWL<20041> A_IWL<20040> A_IWL<20039> A_IWL<20038> A_IWL<20037> A_IWL<20036> A_IWL<20035> A_IWL<20034> A_IWL<20033> A_IWL<20032> A_IWL<20031> A_IWL<20030> A_IWL<20029> A_IWL<20028> A_IWL<20027> A_IWL<20026> A_IWL<20025> A_IWL<20024> A_IWL<20023> A_IWL<20022> A_IWL<20021> A_IWL<20020> A_IWL<20019> A_IWL<20018> A_IWL<20017> A_IWL<20016> A_IWL<20015> A_IWL<20014> A_IWL<20013> A_IWL<20012> A_IWL<20011> A_IWL<20010> A_IWL<20009> A_IWL<20008> A_IWL<20007> A_IWL<20006> A_IWL<20005> A_IWL<20004> A_IWL<20003> A_IWL<20002> A_IWL<20001> A_IWL<20000> A_IWL<19999> A_IWL<19998> A_IWL<19997> A_IWL<19996> A_IWL<19995> A_IWL<19994> A_IWL<19993> A_IWL<19992> A_IWL<19991> A_IWL<19990> A_IWL<19989> A_IWL<19988> A_IWL<19987> A_IWL<19986> A_IWL<19985> A_IWL<19984> A_IWL<19983> A_IWL<19982> A_IWL<19981> A_IWL<19980> A_IWL<19979> A_IWL<19978> A_IWL<19977> A_IWL<19976> A_IWL<19975> A_IWL<19974> A_IWL<19973> A_IWL<19972> A_IWL<19971> A_IWL<19970> A_IWL<19969> A_IWL<19968> A_IWL<20991> A_IWL<20990> A_IWL<20989> A_IWL<20988> A_IWL<20987> A_IWL<20986> A_IWL<20985> A_IWL<20984> A_IWL<20983> A_IWL<20982> A_IWL<20981> A_IWL<20980> A_IWL<20979> A_IWL<20978> A_IWL<20977> A_IWL<20976> A_IWL<20975> A_IWL<20974> A_IWL<20973> A_IWL<20972> A_IWL<20971> A_IWL<20970> A_IWL<20969> A_IWL<20968> A_IWL<20967> A_IWL<20966> A_IWL<20965> A_IWL<20964> A_IWL<20963> A_IWL<20962> A_IWL<20961> A_IWL<20960> A_IWL<20959> A_IWL<20958> A_IWL<20957> A_IWL<20956> A_IWL<20955> A_IWL<20954> A_IWL<20953> A_IWL<20952> A_IWL<20951> A_IWL<20950> A_IWL<20949> A_IWL<20948> A_IWL<20947> A_IWL<20946> A_IWL<20945> A_IWL<20944> A_IWL<20943> A_IWL<20942> A_IWL<20941> A_IWL<20940> A_IWL<20939> A_IWL<20938> A_IWL<20937> A_IWL<20936> A_IWL<20935> A_IWL<20934> A_IWL<20933> A_IWL<20932> A_IWL<20931> A_IWL<20930> A_IWL<20929> A_IWL<20928> A_IWL<20927> A_IWL<20926> A_IWL<20925> A_IWL<20924> A_IWL<20923> A_IWL<20922> A_IWL<20921> A_IWL<20920> A_IWL<20919> A_IWL<20918> A_IWL<20917> A_IWL<20916> A_IWL<20915> A_IWL<20914> A_IWL<20913> A_IWL<20912> A_IWL<20911> A_IWL<20910> A_IWL<20909> A_IWL<20908> A_IWL<20907> A_IWL<20906> A_IWL<20905> A_IWL<20904> A_IWL<20903> A_IWL<20902> A_IWL<20901> A_IWL<20900> A_IWL<20899> A_IWL<20898> A_IWL<20897> A_IWL<20896> A_IWL<20895> A_IWL<20894> A_IWL<20893> A_IWL<20892> A_IWL<20891> A_IWL<20890> A_IWL<20889> A_IWL<20888> A_IWL<20887> A_IWL<20886> A_IWL<20885> A_IWL<20884> A_IWL<20883> A_IWL<20882> A_IWL<20881> A_IWL<20880> A_IWL<20879> A_IWL<20878> A_IWL<20877> A_IWL<20876> A_IWL<20875> A_IWL<20874> A_IWL<20873> A_IWL<20872> A_IWL<20871> A_IWL<20870> A_IWL<20869> A_IWL<20868> A_IWL<20867> A_IWL<20866> A_IWL<20865> A_IWL<20864> A_IWL<20863> A_IWL<20862> A_IWL<20861> A_IWL<20860> A_IWL<20859> A_IWL<20858> A_IWL<20857> A_IWL<20856> A_IWL<20855> A_IWL<20854> A_IWL<20853> A_IWL<20852> A_IWL<20851> A_IWL<20850> A_IWL<20849> A_IWL<20848> A_IWL<20847> A_IWL<20846> A_IWL<20845> A_IWL<20844> A_IWL<20843> A_IWL<20842> A_IWL<20841> A_IWL<20840> A_IWL<20839> A_IWL<20838> A_IWL<20837> A_IWL<20836> A_IWL<20835> A_IWL<20834> A_IWL<20833> A_IWL<20832> A_IWL<20831> A_IWL<20830> A_IWL<20829> A_IWL<20828> A_IWL<20827> A_IWL<20826> A_IWL<20825> A_IWL<20824> A_IWL<20823> A_IWL<20822> A_IWL<20821> A_IWL<20820> A_IWL<20819> A_IWL<20818> A_IWL<20817> A_IWL<20816> A_IWL<20815> A_IWL<20814> A_IWL<20813> A_IWL<20812> A_IWL<20811> A_IWL<20810> A_IWL<20809> A_IWL<20808> A_IWL<20807> A_IWL<20806> A_IWL<20805> A_IWL<20804> A_IWL<20803> A_IWL<20802> A_IWL<20801> A_IWL<20800> A_IWL<20799> A_IWL<20798> A_IWL<20797> A_IWL<20796> A_IWL<20795> A_IWL<20794> A_IWL<20793> A_IWL<20792> A_IWL<20791> A_IWL<20790> A_IWL<20789> A_IWL<20788> A_IWL<20787> A_IWL<20786> A_IWL<20785> A_IWL<20784> A_IWL<20783> A_IWL<20782> A_IWL<20781> A_IWL<20780> A_IWL<20779> A_IWL<20778> A_IWL<20777> A_IWL<20776> A_IWL<20775> A_IWL<20774> A_IWL<20773> A_IWL<20772> A_IWL<20771> A_IWL<20770> A_IWL<20769> A_IWL<20768> A_IWL<20767> A_IWL<20766> A_IWL<20765> A_IWL<20764> A_IWL<20763> A_IWL<20762> A_IWL<20761> A_IWL<20760> A_IWL<20759> A_IWL<20758> A_IWL<20757> A_IWL<20756> A_IWL<20755> A_IWL<20754> A_IWL<20753> A_IWL<20752> A_IWL<20751> A_IWL<20750> A_IWL<20749> A_IWL<20748> A_IWL<20747> A_IWL<20746> A_IWL<20745> A_IWL<20744> A_IWL<20743> A_IWL<20742> A_IWL<20741> A_IWL<20740> A_IWL<20739> A_IWL<20738> A_IWL<20737> A_IWL<20736> A_IWL<20735> A_IWL<20734> A_IWL<20733> A_IWL<20732> A_IWL<20731> A_IWL<20730> A_IWL<20729> A_IWL<20728> A_IWL<20727> A_IWL<20726> A_IWL<20725> A_IWL<20724> A_IWL<20723> A_IWL<20722> A_IWL<20721> A_IWL<20720> A_IWL<20719> A_IWL<20718> A_IWL<20717> A_IWL<20716> A_IWL<20715> A_IWL<20714> A_IWL<20713> A_IWL<20712> A_IWL<20711> A_IWL<20710> A_IWL<20709> A_IWL<20708> A_IWL<20707> A_IWL<20706> A_IWL<20705> A_IWL<20704> A_IWL<20703> A_IWL<20702> A_IWL<20701> A_IWL<20700> A_IWL<20699> A_IWL<20698> A_IWL<20697> A_IWL<20696> A_IWL<20695> A_IWL<20694> A_IWL<20693> A_IWL<20692> A_IWL<20691> A_IWL<20690> A_IWL<20689> A_IWL<20688> A_IWL<20687> A_IWL<20686> A_IWL<20685> A_IWL<20684> A_IWL<20683> A_IWL<20682> A_IWL<20681> A_IWL<20680> A_IWL<20679> A_IWL<20678> A_IWL<20677> A_IWL<20676> A_IWL<20675> A_IWL<20674> A_IWL<20673> A_IWL<20672> A_IWL<20671> A_IWL<20670> A_IWL<20669> A_IWL<20668> A_IWL<20667> A_IWL<20666> A_IWL<20665> A_IWL<20664> A_IWL<20663> A_IWL<20662> A_IWL<20661> A_IWL<20660> A_IWL<20659> A_IWL<20658> A_IWL<20657> A_IWL<20656> A_IWL<20655> A_IWL<20654> A_IWL<20653> A_IWL<20652> A_IWL<20651> A_IWL<20650> A_IWL<20649> A_IWL<20648> A_IWL<20647> A_IWL<20646> A_IWL<20645> A_IWL<20644> A_IWL<20643> A_IWL<20642> A_IWL<20641> A_IWL<20640> A_IWL<20639> A_IWL<20638> A_IWL<20637> A_IWL<20636> A_IWL<20635> A_IWL<20634> A_IWL<20633> A_IWL<20632> A_IWL<20631> A_IWL<20630> A_IWL<20629> A_IWL<20628> A_IWL<20627> A_IWL<20626> A_IWL<20625> A_IWL<20624> A_IWL<20623> A_IWL<20622> A_IWL<20621> A_IWL<20620> A_IWL<20619> A_IWL<20618> A_IWL<20617> A_IWL<20616> A_IWL<20615> A_IWL<20614> A_IWL<20613> A_IWL<20612> A_IWL<20611> A_IWL<20610> A_IWL<20609> A_IWL<20608> A_IWL<20607> A_IWL<20606> A_IWL<20605> A_IWL<20604> A_IWL<20603> A_IWL<20602> A_IWL<20601> A_IWL<20600> A_IWL<20599> A_IWL<20598> A_IWL<20597> A_IWL<20596> A_IWL<20595> A_IWL<20594> A_IWL<20593> A_IWL<20592> A_IWL<20591> A_IWL<20590> A_IWL<20589> A_IWL<20588> A_IWL<20587> A_IWL<20586> A_IWL<20585> A_IWL<20584> A_IWL<20583> A_IWL<20582> A_IWL<20581> A_IWL<20580> A_IWL<20579> A_IWL<20578> A_IWL<20577> A_IWL<20576> A_IWL<20575> A_IWL<20574> A_IWL<20573> A_IWL<20572> A_IWL<20571> A_IWL<20570> A_IWL<20569> A_IWL<20568> A_IWL<20567> A_IWL<20566> A_IWL<20565> A_IWL<20564> A_IWL<20563> A_IWL<20562> A_IWL<20561> A_IWL<20560> A_IWL<20559> A_IWL<20558> A_IWL<20557> A_IWL<20556> A_IWL<20555> A_IWL<20554> A_IWL<20553> A_IWL<20552> A_IWL<20551> A_IWL<20550> A_IWL<20549> A_IWL<20548> A_IWL<20547> A_IWL<20546> A_IWL<20545> A_IWL<20544> A_IWL<20543> A_IWL<20542> A_IWL<20541> A_IWL<20540> A_IWL<20539> A_IWL<20538> A_IWL<20537> A_IWL<20536> A_IWL<20535> A_IWL<20534> A_IWL<20533> A_IWL<20532> A_IWL<20531> A_IWL<20530> A_IWL<20529> A_IWL<20528> A_IWL<20527> A_IWL<20526> A_IWL<20525> A_IWL<20524> A_IWL<20523> A_IWL<20522> A_IWL<20521> A_IWL<20520> A_IWL<20519> A_IWL<20518> A_IWL<20517> A_IWL<20516> A_IWL<20515> A_IWL<20514> A_IWL<20513> A_IWL<20512> A_IWL<20511> A_IWL<20510> A_IWL<20509> A_IWL<20508> A_IWL<20507> A_IWL<20506> A_IWL<20505> A_IWL<20504> A_IWL<20503> A_IWL<20502> A_IWL<20501> A_IWL<20500> A_IWL<20499> A_IWL<20498> A_IWL<20497> A_IWL<20496> A_IWL<20495> A_IWL<20494> A_IWL<20493> A_IWL<20492> A_IWL<20491> A_IWL<20490> A_IWL<20489> A_IWL<20488> A_IWL<20487> A_IWL<20486> A_IWL<20485> A_IWL<20484> A_IWL<20483> A_IWL<20482> A_IWL<20481> A_IWL<20480> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<39> A_BLC<79> A_BLC<78> A_BLC_TOP<79> A_BLC_TOP<78> A_BLT<79> A_BLT<78> A_BLT_TOP<79> A_BLT_TOP<78> A_IWL<19967> A_IWL<19966> A_IWL<19965> A_IWL<19964> A_IWL<19963> A_IWL<19962> A_IWL<19961> A_IWL<19960> A_IWL<19959> A_IWL<19958> A_IWL<19957> A_IWL<19956> A_IWL<19955> A_IWL<19954> A_IWL<19953> A_IWL<19952> A_IWL<19951> A_IWL<19950> A_IWL<19949> A_IWL<19948> A_IWL<19947> A_IWL<19946> A_IWL<19945> A_IWL<19944> A_IWL<19943> A_IWL<19942> A_IWL<19941> A_IWL<19940> A_IWL<19939> A_IWL<19938> A_IWL<19937> A_IWL<19936> A_IWL<19935> A_IWL<19934> A_IWL<19933> A_IWL<19932> A_IWL<19931> A_IWL<19930> A_IWL<19929> A_IWL<19928> A_IWL<19927> A_IWL<19926> A_IWL<19925> A_IWL<19924> A_IWL<19923> A_IWL<19922> A_IWL<19921> A_IWL<19920> A_IWL<19919> A_IWL<19918> A_IWL<19917> A_IWL<19916> A_IWL<19915> A_IWL<19914> A_IWL<19913> A_IWL<19912> A_IWL<19911> A_IWL<19910> A_IWL<19909> A_IWL<19908> A_IWL<19907> A_IWL<19906> A_IWL<19905> A_IWL<19904> A_IWL<19903> A_IWL<19902> A_IWL<19901> A_IWL<19900> A_IWL<19899> A_IWL<19898> A_IWL<19897> A_IWL<19896> A_IWL<19895> A_IWL<19894> A_IWL<19893> A_IWL<19892> A_IWL<19891> A_IWL<19890> A_IWL<19889> A_IWL<19888> A_IWL<19887> A_IWL<19886> A_IWL<19885> A_IWL<19884> A_IWL<19883> A_IWL<19882> A_IWL<19881> A_IWL<19880> A_IWL<19879> A_IWL<19878> A_IWL<19877> A_IWL<19876> A_IWL<19875> A_IWL<19874> A_IWL<19873> A_IWL<19872> A_IWL<19871> A_IWL<19870> A_IWL<19869> A_IWL<19868> A_IWL<19867> A_IWL<19866> A_IWL<19865> A_IWL<19864> A_IWL<19863> A_IWL<19862> A_IWL<19861> A_IWL<19860> A_IWL<19859> A_IWL<19858> A_IWL<19857> A_IWL<19856> A_IWL<19855> A_IWL<19854> A_IWL<19853> A_IWL<19852> A_IWL<19851> A_IWL<19850> A_IWL<19849> A_IWL<19848> A_IWL<19847> A_IWL<19846> A_IWL<19845> A_IWL<19844> A_IWL<19843> A_IWL<19842> A_IWL<19841> A_IWL<19840> A_IWL<19839> A_IWL<19838> A_IWL<19837> A_IWL<19836> A_IWL<19835> A_IWL<19834> A_IWL<19833> A_IWL<19832> A_IWL<19831> A_IWL<19830> A_IWL<19829> A_IWL<19828> A_IWL<19827> A_IWL<19826> A_IWL<19825> A_IWL<19824> A_IWL<19823> A_IWL<19822> A_IWL<19821> A_IWL<19820> A_IWL<19819> A_IWL<19818> A_IWL<19817> A_IWL<19816> A_IWL<19815> A_IWL<19814> A_IWL<19813> A_IWL<19812> A_IWL<19811> A_IWL<19810> A_IWL<19809> A_IWL<19808> A_IWL<19807> A_IWL<19806> A_IWL<19805> A_IWL<19804> A_IWL<19803> A_IWL<19802> A_IWL<19801> A_IWL<19800> A_IWL<19799> A_IWL<19798> A_IWL<19797> A_IWL<19796> A_IWL<19795> A_IWL<19794> A_IWL<19793> A_IWL<19792> A_IWL<19791> A_IWL<19790> A_IWL<19789> A_IWL<19788> A_IWL<19787> A_IWL<19786> A_IWL<19785> A_IWL<19784> A_IWL<19783> A_IWL<19782> A_IWL<19781> A_IWL<19780> A_IWL<19779> A_IWL<19778> A_IWL<19777> A_IWL<19776> A_IWL<19775> A_IWL<19774> A_IWL<19773> A_IWL<19772> A_IWL<19771> A_IWL<19770> A_IWL<19769> A_IWL<19768> A_IWL<19767> A_IWL<19766> A_IWL<19765> A_IWL<19764> A_IWL<19763> A_IWL<19762> A_IWL<19761> A_IWL<19760> A_IWL<19759> A_IWL<19758> A_IWL<19757> A_IWL<19756> A_IWL<19755> A_IWL<19754> A_IWL<19753> A_IWL<19752> A_IWL<19751> A_IWL<19750> A_IWL<19749> A_IWL<19748> A_IWL<19747> A_IWL<19746> A_IWL<19745> A_IWL<19744> A_IWL<19743> A_IWL<19742> A_IWL<19741> A_IWL<19740> A_IWL<19739> A_IWL<19738> A_IWL<19737> A_IWL<19736> A_IWL<19735> A_IWL<19734> A_IWL<19733> A_IWL<19732> A_IWL<19731> A_IWL<19730> A_IWL<19729> A_IWL<19728> A_IWL<19727> A_IWL<19726> A_IWL<19725> A_IWL<19724> A_IWL<19723> A_IWL<19722> A_IWL<19721> A_IWL<19720> A_IWL<19719> A_IWL<19718> A_IWL<19717> A_IWL<19716> A_IWL<19715> A_IWL<19714> A_IWL<19713> A_IWL<19712> A_IWL<19711> A_IWL<19710> A_IWL<19709> A_IWL<19708> A_IWL<19707> A_IWL<19706> A_IWL<19705> A_IWL<19704> A_IWL<19703> A_IWL<19702> A_IWL<19701> A_IWL<19700> A_IWL<19699> A_IWL<19698> A_IWL<19697> A_IWL<19696> A_IWL<19695> A_IWL<19694> A_IWL<19693> A_IWL<19692> A_IWL<19691> A_IWL<19690> A_IWL<19689> A_IWL<19688> A_IWL<19687> A_IWL<19686> A_IWL<19685> A_IWL<19684> A_IWL<19683> A_IWL<19682> A_IWL<19681> A_IWL<19680> A_IWL<19679> A_IWL<19678> A_IWL<19677> A_IWL<19676> A_IWL<19675> A_IWL<19674> A_IWL<19673> A_IWL<19672> A_IWL<19671> A_IWL<19670> A_IWL<19669> A_IWL<19668> A_IWL<19667> A_IWL<19666> A_IWL<19665> A_IWL<19664> A_IWL<19663> A_IWL<19662> A_IWL<19661> A_IWL<19660> A_IWL<19659> A_IWL<19658> A_IWL<19657> A_IWL<19656> A_IWL<19655> A_IWL<19654> A_IWL<19653> A_IWL<19652> A_IWL<19651> A_IWL<19650> A_IWL<19649> A_IWL<19648> A_IWL<19647> A_IWL<19646> A_IWL<19645> A_IWL<19644> A_IWL<19643> A_IWL<19642> A_IWL<19641> A_IWL<19640> A_IWL<19639> A_IWL<19638> A_IWL<19637> A_IWL<19636> A_IWL<19635> A_IWL<19634> A_IWL<19633> A_IWL<19632> A_IWL<19631> A_IWL<19630> A_IWL<19629> A_IWL<19628> A_IWL<19627> A_IWL<19626> A_IWL<19625> A_IWL<19624> A_IWL<19623> A_IWL<19622> A_IWL<19621> A_IWL<19620> A_IWL<19619> A_IWL<19618> A_IWL<19617> A_IWL<19616> A_IWL<19615> A_IWL<19614> A_IWL<19613> A_IWL<19612> A_IWL<19611> A_IWL<19610> A_IWL<19609> A_IWL<19608> A_IWL<19607> A_IWL<19606> A_IWL<19605> A_IWL<19604> A_IWL<19603> A_IWL<19602> A_IWL<19601> A_IWL<19600> A_IWL<19599> A_IWL<19598> A_IWL<19597> A_IWL<19596> A_IWL<19595> A_IWL<19594> A_IWL<19593> A_IWL<19592> A_IWL<19591> A_IWL<19590> A_IWL<19589> A_IWL<19588> A_IWL<19587> A_IWL<19586> A_IWL<19585> A_IWL<19584> A_IWL<19583> A_IWL<19582> A_IWL<19581> A_IWL<19580> A_IWL<19579> A_IWL<19578> A_IWL<19577> A_IWL<19576> A_IWL<19575> A_IWL<19574> A_IWL<19573> A_IWL<19572> A_IWL<19571> A_IWL<19570> A_IWL<19569> A_IWL<19568> A_IWL<19567> A_IWL<19566> A_IWL<19565> A_IWL<19564> A_IWL<19563> A_IWL<19562> A_IWL<19561> A_IWL<19560> A_IWL<19559> A_IWL<19558> A_IWL<19557> A_IWL<19556> A_IWL<19555> A_IWL<19554> A_IWL<19553> A_IWL<19552> A_IWL<19551> A_IWL<19550> A_IWL<19549> A_IWL<19548> A_IWL<19547> A_IWL<19546> A_IWL<19545> A_IWL<19544> A_IWL<19543> A_IWL<19542> A_IWL<19541> A_IWL<19540> A_IWL<19539> A_IWL<19538> A_IWL<19537> A_IWL<19536> A_IWL<19535> A_IWL<19534> A_IWL<19533> A_IWL<19532> A_IWL<19531> A_IWL<19530> A_IWL<19529> A_IWL<19528> A_IWL<19527> A_IWL<19526> A_IWL<19525> A_IWL<19524> A_IWL<19523> A_IWL<19522> A_IWL<19521> A_IWL<19520> A_IWL<19519> A_IWL<19518> A_IWL<19517> A_IWL<19516> A_IWL<19515> A_IWL<19514> A_IWL<19513> A_IWL<19512> A_IWL<19511> A_IWL<19510> A_IWL<19509> A_IWL<19508> A_IWL<19507> A_IWL<19506> A_IWL<19505> A_IWL<19504> A_IWL<19503> A_IWL<19502> A_IWL<19501> A_IWL<19500> A_IWL<19499> A_IWL<19498> A_IWL<19497> A_IWL<19496> A_IWL<19495> A_IWL<19494> A_IWL<19493> A_IWL<19492> A_IWL<19491> A_IWL<19490> A_IWL<19489> A_IWL<19488> A_IWL<19487> A_IWL<19486> A_IWL<19485> A_IWL<19484> A_IWL<19483> A_IWL<19482> A_IWL<19481> A_IWL<19480> A_IWL<19479> A_IWL<19478> A_IWL<19477> A_IWL<19476> A_IWL<19475> A_IWL<19474> A_IWL<19473> A_IWL<19472> A_IWL<19471> A_IWL<19470> A_IWL<19469> A_IWL<19468> A_IWL<19467> A_IWL<19466> A_IWL<19465> A_IWL<19464> A_IWL<19463> A_IWL<19462> A_IWL<19461> A_IWL<19460> A_IWL<19459> A_IWL<19458> A_IWL<19457> A_IWL<19456> A_IWL<20479> A_IWL<20478> A_IWL<20477> A_IWL<20476> A_IWL<20475> A_IWL<20474> A_IWL<20473> A_IWL<20472> A_IWL<20471> A_IWL<20470> A_IWL<20469> A_IWL<20468> A_IWL<20467> A_IWL<20466> A_IWL<20465> A_IWL<20464> A_IWL<20463> A_IWL<20462> A_IWL<20461> A_IWL<20460> A_IWL<20459> A_IWL<20458> A_IWL<20457> A_IWL<20456> A_IWL<20455> A_IWL<20454> A_IWL<20453> A_IWL<20452> A_IWL<20451> A_IWL<20450> A_IWL<20449> A_IWL<20448> A_IWL<20447> A_IWL<20446> A_IWL<20445> A_IWL<20444> A_IWL<20443> A_IWL<20442> A_IWL<20441> A_IWL<20440> A_IWL<20439> A_IWL<20438> A_IWL<20437> A_IWL<20436> A_IWL<20435> A_IWL<20434> A_IWL<20433> A_IWL<20432> A_IWL<20431> A_IWL<20430> A_IWL<20429> A_IWL<20428> A_IWL<20427> A_IWL<20426> A_IWL<20425> A_IWL<20424> A_IWL<20423> A_IWL<20422> A_IWL<20421> A_IWL<20420> A_IWL<20419> A_IWL<20418> A_IWL<20417> A_IWL<20416> A_IWL<20415> A_IWL<20414> A_IWL<20413> A_IWL<20412> A_IWL<20411> A_IWL<20410> A_IWL<20409> A_IWL<20408> A_IWL<20407> A_IWL<20406> A_IWL<20405> A_IWL<20404> A_IWL<20403> A_IWL<20402> A_IWL<20401> A_IWL<20400> A_IWL<20399> A_IWL<20398> A_IWL<20397> A_IWL<20396> A_IWL<20395> A_IWL<20394> A_IWL<20393> A_IWL<20392> A_IWL<20391> A_IWL<20390> A_IWL<20389> A_IWL<20388> A_IWL<20387> A_IWL<20386> A_IWL<20385> A_IWL<20384> A_IWL<20383> A_IWL<20382> A_IWL<20381> A_IWL<20380> A_IWL<20379> A_IWL<20378> A_IWL<20377> A_IWL<20376> A_IWL<20375> A_IWL<20374> A_IWL<20373> A_IWL<20372> A_IWL<20371> A_IWL<20370> A_IWL<20369> A_IWL<20368> A_IWL<20367> A_IWL<20366> A_IWL<20365> A_IWL<20364> A_IWL<20363> A_IWL<20362> A_IWL<20361> A_IWL<20360> A_IWL<20359> A_IWL<20358> A_IWL<20357> A_IWL<20356> A_IWL<20355> A_IWL<20354> A_IWL<20353> A_IWL<20352> A_IWL<20351> A_IWL<20350> A_IWL<20349> A_IWL<20348> A_IWL<20347> A_IWL<20346> A_IWL<20345> A_IWL<20344> A_IWL<20343> A_IWL<20342> A_IWL<20341> A_IWL<20340> A_IWL<20339> A_IWL<20338> A_IWL<20337> A_IWL<20336> A_IWL<20335> A_IWL<20334> A_IWL<20333> A_IWL<20332> A_IWL<20331> A_IWL<20330> A_IWL<20329> A_IWL<20328> A_IWL<20327> A_IWL<20326> A_IWL<20325> A_IWL<20324> A_IWL<20323> A_IWL<20322> A_IWL<20321> A_IWL<20320> A_IWL<20319> A_IWL<20318> A_IWL<20317> A_IWL<20316> A_IWL<20315> A_IWL<20314> A_IWL<20313> A_IWL<20312> A_IWL<20311> A_IWL<20310> A_IWL<20309> A_IWL<20308> A_IWL<20307> A_IWL<20306> A_IWL<20305> A_IWL<20304> A_IWL<20303> A_IWL<20302> A_IWL<20301> A_IWL<20300> A_IWL<20299> A_IWL<20298> A_IWL<20297> A_IWL<20296> A_IWL<20295> A_IWL<20294> A_IWL<20293> A_IWL<20292> A_IWL<20291> A_IWL<20290> A_IWL<20289> A_IWL<20288> A_IWL<20287> A_IWL<20286> A_IWL<20285> A_IWL<20284> A_IWL<20283> A_IWL<20282> A_IWL<20281> A_IWL<20280> A_IWL<20279> A_IWL<20278> A_IWL<20277> A_IWL<20276> A_IWL<20275> A_IWL<20274> A_IWL<20273> A_IWL<20272> A_IWL<20271> A_IWL<20270> A_IWL<20269> A_IWL<20268> A_IWL<20267> A_IWL<20266> A_IWL<20265> A_IWL<20264> A_IWL<20263> A_IWL<20262> A_IWL<20261> A_IWL<20260> A_IWL<20259> A_IWL<20258> A_IWL<20257> A_IWL<20256> A_IWL<20255> A_IWL<20254> A_IWL<20253> A_IWL<20252> A_IWL<20251> A_IWL<20250> A_IWL<20249> A_IWL<20248> A_IWL<20247> A_IWL<20246> A_IWL<20245> A_IWL<20244> A_IWL<20243> A_IWL<20242> A_IWL<20241> A_IWL<20240> A_IWL<20239> A_IWL<20238> A_IWL<20237> A_IWL<20236> A_IWL<20235> A_IWL<20234> A_IWL<20233> A_IWL<20232> A_IWL<20231> A_IWL<20230> A_IWL<20229> A_IWL<20228> A_IWL<20227> A_IWL<20226> A_IWL<20225> A_IWL<20224> A_IWL<20223> A_IWL<20222> A_IWL<20221> A_IWL<20220> A_IWL<20219> A_IWL<20218> A_IWL<20217> A_IWL<20216> A_IWL<20215> A_IWL<20214> A_IWL<20213> A_IWL<20212> A_IWL<20211> A_IWL<20210> A_IWL<20209> A_IWL<20208> A_IWL<20207> A_IWL<20206> A_IWL<20205> A_IWL<20204> A_IWL<20203> A_IWL<20202> A_IWL<20201> A_IWL<20200> A_IWL<20199> A_IWL<20198> A_IWL<20197> A_IWL<20196> A_IWL<20195> A_IWL<20194> A_IWL<20193> A_IWL<20192> A_IWL<20191> A_IWL<20190> A_IWL<20189> A_IWL<20188> A_IWL<20187> A_IWL<20186> A_IWL<20185> A_IWL<20184> A_IWL<20183> A_IWL<20182> A_IWL<20181> A_IWL<20180> A_IWL<20179> A_IWL<20178> A_IWL<20177> A_IWL<20176> A_IWL<20175> A_IWL<20174> A_IWL<20173> A_IWL<20172> A_IWL<20171> A_IWL<20170> A_IWL<20169> A_IWL<20168> A_IWL<20167> A_IWL<20166> A_IWL<20165> A_IWL<20164> A_IWL<20163> A_IWL<20162> A_IWL<20161> A_IWL<20160> A_IWL<20159> A_IWL<20158> A_IWL<20157> A_IWL<20156> A_IWL<20155> A_IWL<20154> A_IWL<20153> A_IWL<20152> A_IWL<20151> A_IWL<20150> A_IWL<20149> A_IWL<20148> A_IWL<20147> A_IWL<20146> A_IWL<20145> A_IWL<20144> A_IWL<20143> A_IWL<20142> A_IWL<20141> A_IWL<20140> A_IWL<20139> A_IWL<20138> A_IWL<20137> A_IWL<20136> A_IWL<20135> A_IWL<20134> A_IWL<20133> A_IWL<20132> A_IWL<20131> A_IWL<20130> A_IWL<20129> A_IWL<20128> A_IWL<20127> A_IWL<20126> A_IWL<20125> A_IWL<20124> A_IWL<20123> A_IWL<20122> A_IWL<20121> A_IWL<20120> A_IWL<20119> A_IWL<20118> A_IWL<20117> A_IWL<20116> A_IWL<20115> A_IWL<20114> A_IWL<20113> A_IWL<20112> A_IWL<20111> A_IWL<20110> A_IWL<20109> A_IWL<20108> A_IWL<20107> A_IWL<20106> A_IWL<20105> A_IWL<20104> A_IWL<20103> A_IWL<20102> A_IWL<20101> A_IWL<20100> A_IWL<20099> A_IWL<20098> A_IWL<20097> A_IWL<20096> A_IWL<20095> A_IWL<20094> A_IWL<20093> A_IWL<20092> A_IWL<20091> A_IWL<20090> A_IWL<20089> A_IWL<20088> A_IWL<20087> A_IWL<20086> A_IWL<20085> A_IWL<20084> A_IWL<20083> A_IWL<20082> A_IWL<20081> A_IWL<20080> A_IWL<20079> A_IWL<20078> A_IWL<20077> A_IWL<20076> A_IWL<20075> A_IWL<20074> A_IWL<20073> A_IWL<20072> A_IWL<20071> A_IWL<20070> A_IWL<20069> A_IWL<20068> A_IWL<20067> A_IWL<20066> A_IWL<20065> A_IWL<20064> A_IWL<20063> A_IWL<20062> A_IWL<20061> A_IWL<20060> A_IWL<20059> A_IWL<20058> A_IWL<20057> A_IWL<20056> A_IWL<20055> A_IWL<20054> A_IWL<20053> A_IWL<20052> A_IWL<20051> A_IWL<20050> A_IWL<20049> A_IWL<20048> A_IWL<20047> A_IWL<20046> A_IWL<20045> A_IWL<20044> A_IWL<20043> A_IWL<20042> A_IWL<20041> A_IWL<20040> A_IWL<20039> A_IWL<20038> A_IWL<20037> A_IWL<20036> A_IWL<20035> A_IWL<20034> A_IWL<20033> A_IWL<20032> A_IWL<20031> A_IWL<20030> A_IWL<20029> A_IWL<20028> A_IWL<20027> A_IWL<20026> A_IWL<20025> A_IWL<20024> A_IWL<20023> A_IWL<20022> A_IWL<20021> A_IWL<20020> A_IWL<20019> A_IWL<20018> A_IWL<20017> A_IWL<20016> A_IWL<20015> A_IWL<20014> A_IWL<20013> A_IWL<20012> A_IWL<20011> A_IWL<20010> A_IWL<20009> A_IWL<20008> A_IWL<20007> A_IWL<20006> A_IWL<20005> A_IWL<20004> A_IWL<20003> A_IWL<20002> A_IWL<20001> A_IWL<20000> A_IWL<19999> A_IWL<19998> A_IWL<19997> A_IWL<19996> A_IWL<19995> A_IWL<19994> A_IWL<19993> A_IWL<19992> A_IWL<19991> A_IWL<19990> A_IWL<19989> A_IWL<19988> A_IWL<19987> A_IWL<19986> A_IWL<19985> A_IWL<19984> A_IWL<19983> A_IWL<19982> A_IWL<19981> A_IWL<19980> A_IWL<19979> A_IWL<19978> A_IWL<19977> A_IWL<19976> A_IWL<19975> A_IWL<19974> A_IWL<19973> A_IWL<19972> A_IWL<19971> A_IWL<19970> A_IWL<19969> A_IWL<19968> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<38> A_BLC<77> A_BLC<76> A_BLC_TOP<77> A_BLC_TOP<76> A_BLT<77> A_BLT<76> A_BLT_TOP<77> A_BLT_TOP<76> A_IWL<19455> A_IWL<19454> A_IWL<19453> A_IWL<19452> A_IWL<19451> A_IWL<19450> A_IWL<19449> A_IWL<19448> A_IWL<19447> A_IWL<19446> A_IWL<19445> A_IWL<19444> A_IWL<19443> A_IWL<19442> A_IWL<19441> A_IWL<19440> A_IWL<19439> A_IWL<19438> A_IWL<19437> A_IWL<19436> A_IWL<19435> A_IWL<19434> A_IWL<19433> A_IWL<19432> A_IWL<19431> A_IWL<19430> A_IWL<19429> A_IWL<19428> A_IWL<19427> A_IWL<19426> A_IWL<19425> A_IWL<19424> A_IWL<19423> A_IWL<19422> A_IWL<19421> A_IWL<19420> A_IWL<19419> A_IWL<19418> A_IWL<19417> A_IWL<19416> A_IWL<19415> A_IWL<19414> A_IWL<19413> A_IWL<19412> A_IWL<19411> A_IWL<19410> A_IWL<19409> A_IWL<19408> A_IWL<19407> A_IWL<19406> A_IWL<19405> A_IWL<19404> A_IWL<19403> A_IWL<19402> A_IWL<19401> A_IWL<19400> A_IWL<19399> A_IWL<19398> A_IWL<19397> A_IWL<19396> A_IWL<19395> A_IWL<19394> A_IWL<19393> A_IWL<19392> A_IWL<19391> A_IWL<19390> A_IWL<19389> A_IWL<19388> A_IWL<19387> A_IWL<19386> A_IWL<19385> A_IWL<19384> A_IWL<19383> A_IWL<19382> A_IWL<19381> A_IWL<19380> A_IWL<19379> A_IWL<19378> A_IWL<19377> A_IWL<19376> A_IWL<19375> A_IWL<19374> A_IWL<19373> A_IWL<19372> A_IWL<19371> A_IWL<19370> A_IWL<19369> A_IWL<19368> A_IWL<19367> A_IWL<19366> A_IWL<19365> A_IWL<19364> A_IWL<19363> A_IWL<19362> A_IWL<19361> A_IWL<19360> A_IWL<19359> A_IWL<19358> A_IWL<19357> A_IWL<19356> A_IWL<19355> A_IWL<19354> A_IWL<19353> A_IWL<19352> A_IWL<19351> A_IWL<19350> A_IWL<19349> A_IWL<19348> A_IWL<19347> A_IWL<19346> A_IWL<19345> A_IWL<19344> A_IWL<19343> A_IWL<19342> A_IWL<19341> A_IWL<19340> A_IWL<19339> A_IWL<19338> A_IWL<19337> A_IWL<19336> A_IWL<19335> A_IWL<19334> A_IWL<19333> A_IWL<19332> A_IWL<19331> A_IWL<19330> A_IWL<19329> A_IWL<19328> A_IWL<19327> A_IWL<19326> A_IWL<19325> A_IWL<19324> A_IWL<19323> A_IWL<19322> A_IWL<19321> A_IWL<19320> A_IWL<19319> A_IWL<19318> A_IWL<19317> A_IWL<19316> A_IWL<19315> A_IWL<19314> A_IWL<19313> A_IWL<19312> A_IWL<19311> A_IWL<19310> A_IWL<19309> A_IWL<19308> A_IWL<19307> A_IWL<19306> A_IWL<19305> A_IWL<19304> A_IWL<19303> A_IWL<19302> A_IWL<19301> A_IWL<19300> A_IWL<19299> A_IWL<19298> A_IWL<19297> A_IWL<19296> A_IWL<19295> A_IWL<19294> A_IWL<19293> A_IWL<19292> A_IWL<19291> A_IWL<19290> A_IWL<19289> A_IWL<19288> A_IWL<19287> A_IWL<19286> A_IWL<19285> A_IWL<19284> A_IWL<19283> A_IWL<19282> A_IWL<19281> A_IWL<19280> A_IWL<19279> A_IWL<19278> A_IWL<19277> A_IWL<19276> A_IWL<19275> A_IWL<19274> A_IWL<19273> A_IWL<19272> A_IWL<19271> A_IWL<19270> A_IWL<19269> A_IWL<19268> A_IWL<19267> A_IWL<19266> A_IWL<19265> A_IWL<19264> A_IWL<19263> A_IWL<19262> A_IWL<19261> A_IWL<19260> A_IWL<19259> A_IWL<19258> A_IWL<19257> A_IWL<19256> A_IWL<19255> A_IWL<19254> A_IWL<19253> A_IWL<19252> A_IWL<19251> A_IWL<19250> A_IWL<19249> A_IWL<19248> A_IWL<19247> A_IWL<19246> A_IWL<19245> A_IWL<19244> A_IWL<19243> A_IWL<19242> A_IWL<19241> A_IWL<19240> A_IWL<19239> A_IWL<19238> A_IWL<19237> A_IWL<19236> A_IWL<19235> A_IWL<19234> A_IWL<19233> A_IWL<19232> A_IWL<19231> A_IWL<19230> A_IWL<19229> A_IWL<19228> A_IWL<19227> A_IWL<19226> A_IWL<19225> A_IWL<19224> A_IWL<19223> A_IWL<19222> A_IWL<19221> A_IWL<19220> A_IWL<19219> A_IWL<19218> A_IWL<19217> A_IWL<19216> A_IWL<19215> A_IWL<19214> A_IWL<19213> A_IWL<19212> A_IWL<19211> A_IWL<19210> A_IWL<19209> A_IWL<19208> A_IWL<19207> A_IWL<19206> A_IWL<19205> A_IWL<19204> A_IWL<19203> A_IWL<19202> A_IWL<19201> A_IWL<19200> A_IWL<19199> A_IWL<19198> A_IWL<19197> A_IWL<19196> A_IWL<19195> A_IWL<19194> A_IWL<19193> A_IWL<19192> A_IWL<19191> A_IWL<19190> A_IWL<19189> A_IWL<19188> A_IWL<19187> A_IWL<19186> A_IWL<19185> A_IWL<19184> A_IWL<19183> A_IWL<19182> A_IWL<19181> A_IWL<19180> A_IWL<19179> A_IWL<19178> A_IWL<19177> A_IWL<19176> A_IWL<19175> A_IWL<19174> A_IWL<19173> A_IWL<19172> A_IWL<19171> A_IWL<19170> A_IWL<19169> A_IWL<19168> A_IWL<19167> A_IWL<19166> A_IWL<19165> A_IWL<19164> A_IWL<19163> A_IWL<19162> A_IWL<19161> A_IWL<19160> A_IWL<19159> A_IWL<19158> A_IWL<19157> A_IWL<19156> A_IWL<19155> A_IWL<19154> A_IWL<19153> A_IWL<19152> A_IWL<19151> A_IWL<19150> A_IWL<19149> A_IWL<19148> A_IWL<19147> A_IWL<19146> A_IWL<19145> A_IWL<19144> A_IWL<19143> A_IWL<19142> A_IWL<19141> A_IWL<19140> A_IWL<19139> A_IWL<19138> A_IWL<19137> A_IWL<19136> A_IWL<19135> A_IWL<19134> A_IWL<19133> A_IWL<19132> A_IWL<19131> A_IWL<19130> A_IWL<19129> A_IWL<19128> A_IWL<19127> A_IWL<19126> A_IWL<19125> A_IWL<19124> A_IWL<19123> A_IWL<19122> A_IWL<19121> A_IWL<19120> A_IWL<19119> A_IWL<19118> A_IWL<19117> A_IWL<19116> A_IWL<19115> A_IWL<19114> A_IWL<19113> A_IWL<19112> A_IWL<19111> A_IWL<19110> A_IWL<19109> A_IWL<19108> A_IWL<19107> A_IWL<19106> A_IWL<19105> A_IWL<19104> A_IWL<19103> A_IWL<19102> A_IWL<19101> A_IWL<19100> A_IWL<19099> A_IWL<19098> A_IWL<19097> A_IWL<19096> A_IWL<19095> A_IWL<19094> A_IWL<19093> A_IWL<19092> A_IWL<19091> A_IWL<19090> A_IWL<19089> A_IWL<19088> A_IWL<19087> A_IWL<19086> A_IWL<19085> A_IWL<19084> A_IWL<19083> A_IWL<19082> A_IWL<19081> A_IWL<19080> A_IWL<19079> A_IWL<19078> A_IWL<19077> A_IWL<19076> A_IWL<19075> A_IWL<19074> A_IWL<19073> A_IWL<19072> A_IWL<19071> A_IWL<19070> A_IWL<19069> A_IWL<19068> A_IWL<19067> A_IWL<19066> A_IWL<19065> A_IWL<19064> A_IWL<19063> A_IWL<19062> A_IWL<19061> A_IWL<19060> A_IWL<19059> A_IWL<19058> A_IWL<19057> A_IWL<19056> A_IWL<19055> A_IWL<19054> A_IWL<19053> A_IWL<19052> A_IWL<19051> A_IWL<19050> A_IWL<19049> A_IWL<19048> A_IWL<19047> A_IWL<19046> A_IWL<19045> A_IWL<19044> A_IWL<19043> A_IWL<19042> A_IWL<19041> A_IWL<19040> A_IWL<19039> A_IWL<19038> A_IWL<19037> A_IWL<19036> A_IWL<19035> A_IWL<19034> A_IWL<19033> A_IWL<19032> A_IWL<19031> A_IWL<19030> A_IWL<19029> A_IWL<19028> A_IWL<19027> A_IWL<19026> A_IWL<19025> A_IWL<19024> A_IWL<19023> A_IWL<19022> A_IWL<19021> A_IWL<19020> A_IWL<19019> A_IWL<19018> A_IWL<19017> A_IWL<19016> A_IWL<19015> A_IWL<19014> A_IWL<19013> A_IWL<19012> A_IWL<19011> A_IWL<19010> A_IWL<19009> A_IWL<19008> A_IWL<19007> A_IWL<19006> A_IWL<19005> A_IWL<19004> A_IWL<19003> A_IWL<19002> A_IWL<19001> A_IWL<19000> A_IWL<18999> A_IWL<18998> A_IWL<18997> A_IWL<18996> A_IWL<18995> A_IWL<18994> A_IWL<18993> A_IWL<18992> A_IWL<18991> A_IWL<18990> A_IWL<18989> A_IWL<18988> A_IWL<18987> A_IWL<18986> A_IWL<18985> A_IWL<18984> A_IWL<18983> A_IWL<18982> A_IWL<18981> A_IWL<18980> A_IWL<18979> A_IWL<18978> A_IWL<18977> A_IWL<18976> A_IWL<18975> A_IWL<18974> A_IWL<18973> A_IWL<18972> A_IWL<18971> A_IWL<18970> A_IWL<18969> A_IWL<18968> A_IWL<18967> A_IWL<18966> A_IWL<18965> A_IWL<18964> A_IWL<18963> A_IWL<18962> A_IWL<18961> A_IWL<18960> A_IWL<18959> A_IWL<18958> A_IWL<18957> A_IWL<18956> A_IWL<18955> A_IWL<18954> A_IWL<18953> A_IWL<18952> A_IWL<18951> A_IWL<18950> A_IWL<18949> A_IWL<18948> A_IWL<18947> A_IWL<18946> A_IWL<18945> A_IWL<18944> A_IWL<19967> A_IWL<19966> A_IWL<19965> A_IWL<19964> A_IWL<19963> A_IWL<19962> A_IWL<19961> A_IWL<19960> A_IWL<19959> A_IWL<19958> A_IWL<19957> A_IWL<19956> A_IWL<19955> A_IWL<19954> A_IWL<19953> A_IWL<19952> A_IWL<19951> A_IWL<19950> A_IWL<19949> A_IWL<19948> A_IWL<19947> A_IWL<19946> A_IWL<19945> A_IWL<19944> A_IWL<19943> A_IWL<19942> A_IWL<19941> A_IWL<19940> A_IWL<19939> A_IWL<19938> A_IWL<19937> A_IWL<19936> A_IWL<19935> A_IWL<19934> A_IWL<19933> A_IWL<19932> A_IWL<19931> A_IWL<19930> A_IWL<19929> A_IWL<19928> A_IWL<19927> A_IWL<19926> A_IWL<19925> A_IWL<19924> A_IWL<19923> A_IWL<19922> A_IWL<19921> A_IWL<19920> A_IWL<19919> A_IWL<19918> A_IWL<19917> A_IWL<19916> A_IWL<19915> A_IWL<19914> A_IWL<19913> A_IWL<19912> A_IWL<19911> A_IWL<19910> A_IWL<19909> A_IWL<19908> A_IWL<19907> A_IWL<19906> A_IWL<19905> A_IWL<19904> A_IWL<19903> A_IWL<19902> A_IWL<19901> A_IWL<19900> A_IWL<19899> A_IWL<19898> A_IWL<19897> A_IWL<19896> A_IWL<19895> A_IWL<19894> A_IWL<19893> A_IWL<19892> A_IWL<19891> A_IWL<19890> A_IWL<19889> A_IWL<19888> A_IWL<19887> A_IWL<19886> A_IWL<19885> A_IWL<19884> A_IWL<19883> A_IWL<19882> A_IWL<19881> A_IWL<19880> A_IWL<19879> A_IWL<19878> A_IWL<19877> A_IWL<19876> A_IWL<19875> A_IWL<19874> A_IWL<19873> A_IWL<19872> A_IWL<19871> A_IWL<19870> A_IWL<19869> A_IWL<19868> A_IWL<19867> A_IWL<19866> A_IWL<19865> A_IWL<19864> A_IWL<19863> A_IWL<19862> A_IWL<19861> A_IWL<19860> A_IWL<19859> A_IWL<19858> A_IWL<19857> A_IWL<19856> A_IWL<19855> A_IWL<19854> A_IWL<19853> A_IWL<19852> A_IWL<19851> A_IWL<19850> A_IWL<19849> A_IWL<19848> A_IWL<19847> A_IWL<19846> A_IWL<19845> A_IWL<19844> A_IWL<19843> A_IWL<19842> A_IWL<19841> A_IWL<19840> A_IWL<19839> A_IWL<19838> A_IWL<19837> A_IWL<19836> A_IWL<19835> A_IWL<19834> A_IWL<19833> A_IWL<19832> A_IWL<19831> A_IWL<19830> A_IWL<19829> A_IWL<19828> A_IWL<19827> A_IWL<19826> A_IWL<19825> A_IWL<19824> A_IWL<19823> A_IWL<19822> A_IWL<19821> A_IWL<19820> A_IWL<19819> A_IWL<19818> A_IWL<19817> A_IWL<19816> A_IWL<19815> A_IWL<19814> A_IWL<19813> A_IWL<19812> A_IWL<19811> A_IWL<19810> A_IWL<19809> A_IWL<19808> A_IWL<19807> A_IWL<19806> A_IWL<19805> A_IWL<19804> A_IWL<19803> A_IWL<19802> A_IWL<19801> A_IWL<19800> A_IWL<19799> A_IWL<19798> A_IWL<19797> A_IWL<19796> A_IWL<19795> A_IWL<19794> A_IWL<19793> A_IWL<19792> A_IWL<19791> A_IWL<19790> A_IWL<19789> A_IWL<19788> A_IWL<19787> A_IWL<19786> A_IWL<19785> A_IWL<19784> A_IWL<19783> A_IWL<19782> A_IWL<19781> A_IWL<19780> A_IWL<19779> A_IWL<19778> A_IWL<19777> A_IWL<19776> A_IWL<19775> A_IWL<19774> A_IWL<19773> A_IWL<19772> A_IWL<19771> A_IWL<19770> A_IWL<19769> A_IWL<19768> A_IWL<19767> A_IWL<19766> A_IWL<19765> A_IWL<19764> A_IWL<19763> A_IWL<19762> A_IWL<19761> A_IWL<19760> A_IWL<19759> A_IWL<19758> A_IWL<19757> A_IWL<19756> A_IWL<19755> A_IWL<19754> A_IWL<19753> A_IWL<19752> A_IWL<19751> A_IWL<19750> A_IWL<19749> A_IWL<19748> A_IWL<19747> A_IWL<19746> A_IWL<19745> A_IWL<19744> A_IWL<19743> A_IWL<19742> A_IWL<19741> A_IWL<19740> A_IWL<19739> A_IWL<19738> A_IWL<19737> A_IWL<19736> A_IWL<19735> A_IWL<19734> A_IWL<19733> A_IWL<19732> A_IWL<19731> A_IWL<19730> A_IWL<19729> A_IWL<19728> A_IWL<19727> A_IWL<19726> A_IWL<19725> A_IWL<19724> A_IWL<19723> A_IWL<19722> A_IWL<19721> A_IWL<19720> A_IWL<19719> A_IWL<19718> A_IWL<19717> A_IWL<19716> A_IWL<19715> A_IWL<19714> A_IWL<19713> A_IWL<19712> A_IWL<19711> A_IWL<19710> A_IWL<19709> A_IWL<19708> A_IWL<19707> A_IWL<19706> A_IWL<19705> A_IWL<19704> A_IWL<19703> A_IWL<19702> A_IWL<19701> A_IWL<19700> A_IWL<19699> A_IWL<19698> A_IWL<19697> A_IWL<19696> A_IWL<19695> A_IWL<19694> A_IWL<19693> A_IWL<19692> A_IWL<19691> A_IWL<19690> A_IWL<19689> A_IWL<19688> A_IWL<19687> A_IWL<19686> A_IWL<19685> A_IWL<19684> A_IWL<19683> A_IWL<19682> A_IWL<19681> A_IWL<19680> A_IWL<19679> A_IWL<19678> A_IWL<19677> A_IWL<19676> A_IWL<19675> A_IWL<19674> A_IWL<19673> A_IWL<19672> A_IWL<19671> A_IWL<19670> A_IWL<19669> A_IWL<19668> A_IWL<19667> A_IWL<19666> A_IWL<19665> A_IWL<19664> A_IWL<19663> A_IWL<19662> A_IWL<19661> A_IWL<19660> A_IWL<19659> A_IWL<19658> A_IWL<19657> A_IWL<19656> A_IWL<19655> A_IWL<19654> A_IWL<19653> A_IWL<19652> A_IWL<19651> A_IWL<19650> A_IWL<19649> A_IWL<19648> A_IWL<19647> A_IWL<19646> A_IWL<19645> A_IWL<19644> A_IWL<19643> A_IWL<19642> A_IWL<19641> A_IWL<19640> A_IWL<19639> A_IWL<19638> A_IWL<19637> A_IWL<19636> A_IWL<19635> A_IWL<19634> A_IWL<19633> A_IWL<19632> A_IWL<19631> A_IWL<19630> A_IWL<19629> A_IWL<19628> A_IWL<19627> A_IWL<19626> A_IWL<19625> A_IWL<19624> A_IWL<19623> A_IWL<19622> A_IWL<19621> A_IWL<19620> A_IWL<19619> A_IWL<19618> A_IWL<19617> A_IWL<19616> A_IWL<19615> A_IWL<19614> A_IWL<19613> A_IWL<19612> A_IWL<19611> A_IWL<19610> A_IWL<19609> A_IWL<19608> A_IWL<19607> A_IWL<19606> A_IWL<19605> A_IWL<19604> A_IWL<19603> A_IWL<19602> A_IWL<19601> A_IWL<19600> A_IWL<19599> A_IWL<19598> A_IWL<19597> A_IWL<19596> A_IWL<19595> A_IWL<19594> A_IWL<19593> A_IWL<19592> A_IWL<19591> A_IWL<19590> A_IWL<19589> A_IWL<19588> A_IWL<19587> A_IWL<19586> A_IWL<19585> A_IWL<19584> A_IWL<19583> A_IWL<19582> A_IWL<19581> A_IWL<19580> A_IWL<19579> A_IWL<19578> A_IWL<19577> A_IWL<19576> A_IWL<19575> A_IWL<19574> A_IWL<19573> A_IWL<19572> A_IWL<19571> A_IWL<19570> A_IWL<19569> A_IWL<19568> A_IWL<19567> A_IWL<19566> A_IWL<19565> A_IWL<19564> A_IWL<19563> A_IWL<19562> A_IWL<19561> A_IWL<19560> A_IWL<19559> A_IWL<19558> A_IWL<19557> A_IWL<19556> A_IWL<19555> A_IWL<19554> A_IWL<19553> A_IWL<19552> A_IWL<19551> A_IWL<19550> A_IWL<19549> A_IWL<19548> A_IWL<19547> A_IWL<19546> A_IWL<19545> A_IWL<19544> A_IWL<19543> A_IWL<19542> A_IWL<19541> A_IWL<19540> A_IWL<19539> A_IWL<19538> A_IWL<19537> A_IWL<19536> A_IWL<19535> A_IWL<19534> A_IWL<19533> A_IWL<19532> A_IWL<19531> A_IWL<19530> A_IWL<19529> A_IWL<19528> A_IWL<19527> A_IWL<19526> A_IWL<19525> A_IWL<19524> A_IWL<19523> A_IWL<19522> A_IWL<19521> A_IWL<19520> A_IWL<19519> A_IWL<19518> A_IWL<19517> A_IWL<19516> A_IWL<19515> A_IWL<19514> A_IWL<19513> A_IWL<19512> A_IWL<19511> A_IWL<19510> A_IWL<19509> A_IWL<19508> A_IWL<19507> A_IWL<19506> A_IWL<19505> A_IWL<19504> A_IWL<19503> A_IWL<19502> A_IWL<19501> A_IWL<19500> A_IWL<19499> A_IWL<19498> A_IWL<19497> A_IWL<19496> A_IWL<19495> A_IWL<19494> A_IWL<19493> A_IWL<19492> A_IWL<19491> A_IWL<19490> A_IWL<19489> A_IWL<19488> A_IWL<19487> A_IWL<19486> A_IWL<19485> A_IWL<19484> A_IWL<19483> A_IWL<19482> A_IWL<19481> A_IWL<19480> A_IWL<19479> A_IWL<19478> A_IWL<19477> A_IWL<19476> A_IWL<19475> A_IWL<19474> A_IWL<19473> A_IWL<19472> A_IWL<19471> A_IWL<19470> A_IWL<19469> A_IWL<19468> A_IWL<19467> A_IWL<19466> A_IWL<19465> A_IWL<19464> A_IWL<19463> A_IWL<19462> A_IWL<19461> A_IWL<19460> A_IWL<19459> A_IWL<19458> A_IWL<19457> A_IWL<19456> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<37> A_BLC<75> A_BLC<74> A_BLC_TOP<75> A_BLC_TOP<74> A_BLT<75> A_BLT<74> A_BLT_TOP<75> A_BLT_TOP<74> A_IWL<18943> A_IWL<18942> A_IWL<18941> A_IWL<18940> A_IWL<18939> A_IWL<18938> A_IWL<18937> A_IWL<18936> A_IWL<18935> A_IWL<18934> A_IWL<18933> A_IWL<18932> A_IWL<18931> A_IWL<18930> A_IWL<18929> A_IWL<18928> A_IWL<18927> A_IWL<18926> A_IWL<18925> A_IWL<18924> A_IWL<18923> A_IWL<18922> A_IWL<18921> A_IWL<18920> A_IWL<18919> A_IWL<18918> A_IWL<18917> A_IWL<18916> A_IWL<18915> A_IWL<18914> A_IWL<18913> A_IWL<18912> A_IWL<18911> A_IWL<18910> A_IWL<18909> A_IWL<18908> A_IWL<18907> A_IWL<18906> A_IWL<18905> A_IWL<18904> A_IWL<18903> A_IWL<18902> A_IWL<18901> A_IWL<18900> A_IWL<18899> A_IWL<18898> A_IWL<18897> A_IWL<18896> A_IWL<18895> A_IWL<18894> A_IWL<18893> A_IWL<18892> A_IWL<18891> A_IWL<18890> A_IWL<18889> A_IWL<18888> A_IWL<18887> A_IWL<18886> A_IWL<18885> A_IWL<18884> A_IWL<18883> A_IWL<18882> A_IWL<18881> A_IWL<18880> A_IWL<18879> A_IWL<18878> A_IWL<18877> A_IWL<18876> A_IWL<18875> A_IWL<18874> A_IWL<18873> A_IWL<18872> A_IWL<18871> A_IWL<18870> A_IWL<18869> A_IWL<18868> A_IWL<18867> A_IWL<18866> A_IWL<18865> A_IWL<18864> A_IWL<18863> A_IWL<18862> A_IWL<18861> A_IWL<18860> A_IWL<18859> A_IWL<18858> A_IWL<18857> A_IWL<18856> A_IWL<18855> A_IWL<18854> A_IWL<18853> A_IWL<18852> A_IWL<18851> A_IWL<18850> A_IWL<18849> A_IWL<18848> A_IWL<18847> A_IWL<18846> A_IWL<18845> A_IWL<18844> A_IWL<18843> A_IWL<18842> A_IWL<18841> A_IWL<18840> A_IWL<18839> A_IWL<18838> A_IWL<18837> A_IWL<18836> A_IWL<18835> A_IWL<18834> A_IWL<18833> A_IWL<18832> A_IWL<18831> A_IWL<18830> A_IWL<18829> A_IWL<18828> A_IWL<18827> A_IWL<18826> A_IWL<18825> A_IWL<18824> A_IWL<18823> A_IWL<18822> A_IWL<18821> A_IWL<18820> A_IWL<18819> A_IWL<18818> A_IWL<18817> A_IWL<18816> A_IWL<18815> A_IWL<18814> A_IWL<18813> A_IWL<18812> A_IWL<18811> A_IWL<18810> A_IWL<18809> A_IWL<18808> A_IWL<18807> A_IWL<18806> A_IWL<18805> A_IWL<18804> A_IWL<18803> A_IWL<18802> A_IWL<18801> A_IWL<18800> A_IWL<18799> A_IWL<18798> A_IWL<18797> A_IWL<18796> A_IWL<18795> A_IWL<18794> A_IWL<18793> A_IWL<18792> A_IWL<18791> A_IWL<18790> A_IWL<18789> A_IWL<18788> A_IWL<18787> A_IWL<18786> A_IWL<18785> A_IWL<18784> A_IWL<18783> A_IWL<18782> A_IWL<18781> A_IWL<18780> A_IWL<18779> A_IWL<18778> A_IWL<18777> A_IWL<18776> A_IWL<18775> A_IWL<18774> A_IWL<18773> A_IWL<18772> A_IWL<18771> A_IWL<18770> A_IWL<18769> A_IWL<18768> A_IWL<18767> A_IWL<18766> A_IWL<18765> A_IWL<18764> A_IWL<18763> A_IWL<18762> A_IWL<18761> A_IWL<18760> A_IWL<18759> A_IWL<18758> A_IWL<18757> A_IWL<18756> A_IWL<18755> A_IWL<18754> A_IWL<18753> A_IWL<18752> A_IWL<18751> A_IWL<18750> A_IWL<18749> A_IWL<18748> A_IWL<18747> A_IWL<18746> A_IWL<18745> A_IWL<18744> A_IWL<18743> A_IWL<18742> A_IWL<18741> A_IWL<18740> A_IWL<18739> A_IWL<18738> A_IWL<18737> A_IWL<18736> A_IWL<18735> A_IWL<18734> A_IWL<18733> A_IWL<18732> A_IWL<18731> A_IWL<18730> A_IWL<18729> A_IWL<18728> A_IWL<18727> A_IWL<18726> A_IWL<18725> A_IWL<18724> A_IWL<18723> A_IWL<18722> A_IWL<18721> A_IWL<18720> A_IWL<18719> A_IWL<18718> A_IWL<18717> A_IWL<18716> A_IWL<18715> A_IWL<18714> A_IWL<18713> A_IWL<18712> A_IWL<18711> A_IWL<18710> A_IWL<18709> A_IWL<18708> A_IWL<18707> A_IWL<18706> A_IWL<18705> A_IWL<18704> A_IWL<18703> A_IWL<18702> A_IWL<18701> A_IWL<18700> A_IWL<18699> A_IWL<18698> A_IWL<18697> A_IWL<18696> A_IWL<18695> A_IWL<18694> A_IWL<18693> A_IWL<18692> A_IWL<18691> A_IWL<18690> A_IWL<18689> A_IWL<18688> A_IWL<18687> A_IWL<18686> A_IWL<18685> A_IWL<18684> A_IWL<18683> A_IWL<18682> A_IWL<18681> A_IWL<18680> A_IWL<18679> A_IWL<18678> A_IWL<18677> A_IWL<18676> A_IWL<18675> A_IWL<18674> A_IWL<18673> A_IWL<18672> A_IWL<18671> A_IWL<18670> A_IWL<18669> A_IWL<18668> A_IWL<18667> A_IWL<18666> A_IWL<18665> A_IWL<18664> A_IWL<18663> A_IWL<18662> A_IWL<18661> A_IWL<18660> A_IWL<18659> A_IWL<18658> A_IWL<18657> A_IWL<18656> A_IWL<18655> A_IWL<18654> A_IWL<18653> A_IWL<18652> A_IWL<18651> A_IWL<18650> A_IWL<18649> A_IWL<18648> A_IWL<18647> A_IWL<18646> A_IWL<18645> A_IWL<18644> A_IWL<18643> A_IWL<18642> A_IWL<18641> A_IWL<18640> A_IWL<18639> A_IWL<18638> A_IWL<18637> A_IWL<18636> A_IWL<18635> A_IWL<18634> A_IWL<18633> A_IWL<18632> A_IWL<18631> A_IWL<18630> A_IWL<18629> A_IWL<18628> A_IWL<18627> A_IWL<18626> A_IWL<18625> A_IWL<18624> A_IWL<18623> A_IWL<18622> A_IWL<18621> A_IWL<18620> A_IWL<18619> A_IWL<18618> A_IWL<18617> A_IWL<18616> A_IWL<18615> A_IWL<18614> A_IWL<18613> A_IWL<18612> A_IWL<18611> A_IWL<18610> A_IWL<18609> A_IWL<18608> A_IWL<18607> A_IWL<18606> A_IWL<18605> A_IWL<18604> A_IWL<18603> A_IWL<18602> A_IWL<18601> A_IWL<18600> A_IWL<18599> A_IWL<18598> A_IWL<18597> A_IWL<18596> A_IWL<18595> A_IWL<18594> A_IWL<18593> A_IWL<18592> A_IWL<18591> A_IWL<18590> A_IWL<18589> A_IWL<18588> A_IWL<18587> A_IWL<18586> A_IWL<18585> A_IWL<18584> A_IWL<18583> A_IWL<18582> A_IWL<18581> A_IWL<18580> A_IWL<18579> A_IWL<18578> A_IWL<18577> A_IWL<18576> A_IWL<18575> A_IWL<18574> A_IWL<18573> A_IWL<18572> A_IWL<18571> A_IWL<18570> A_IWL<18569> A_IWL<18568> A_IWL<18567> A_IWL<18566> A_IWL<18565> A_IWL<18564> A_IWL<18563> A_IWL<18562> A_IWL<18561> A_IWL<18560> A_IWL<18559> A_IWL<18558> A_IWL<18557> A_IWL<18556> A_IWL<18555> A_IWL<18554> A_IWL<18553> A_IWL<18552> A_IWL<18551> A_IWL<18550> A_IWL<18549> A_IWL<18548> A_IWL<18547> A_IWL<18546> A_IWL<18545> A_IWL<18544> A_IWL<18543> A_IWL<18542> A_IWL<18541> A_IWL<18540> A_IWL<18539> A_IWL<18538> A_IWL<18537> A_IWL<18536> A_IWL<18535> A_IWL<18534> A_IWL<18533> A_IWL<18532> A_IWL<18531> A_IWL<18530> A_IWL<18529> A_IWL<18528> A_IWL<18527> A_IWL<18526> A_IWL<18525> A_IWL<18524> A_IWL<18523> A_IWL<18522> A_IWL<18521> A_IWL<18520> A_IWL<18519> A_IWL<18518> A_IWL<18517> A_IWL<18516> A_IWL<18515> A_IWL<18514> A_IWL<18513> A_IWL<18512> A_IWL<18511> A_IWL<18510> A_IWL<18509> A_IWL<18508> A_IWL<18507> A_IWL<18506> A_IWL<18505> A_IWL<18504> A_IWL<18503> A_IWL<18502> A_IWL<18501> A_IWL<18500> A_IWL<18499> A_IWL<18498> A_IWL<18497> A_IWL<18496> A_IWL<18495> A_IWL<18494> A_IWL<18493> A_IWL<18492> A_IWL<18491> A_IWL<18490> A_IWL<18489> A_IWL<18488> A_IWL<18487> A_IWL<18486> A_IWL<18485> A_IWL<18484> A_IWL<18483> A_IWL<18482> A_IWL<18481> A_IWL<18480> A_IWL<18479> A_IWL<18478> A_IWL<18477> A_IWL<18476> A_IWL<18475> A_IWL<18474> A_IWL<18473> A_IWL<18472> A_IWL<18471> A_IWL<18470> A_IWL<18469> A_IWL<18468> A_IWL<18467> A_IWL<18466> A_IWL<18465> A_IWL<18464> A_IWL<18463> A_IWL<18462> A_IWL<18461> A_IWL<18460> A_IWL<18459> A_IWL<18458> A_IWL<18457> A_IWL<18456> A_IWL<18455> A_IWL<18454> A_IWL<18453> A_IWL<18452> A_IWL<18451> A_IWL<18450> A_IWL<18449> A_IWL<18448> A_IWL<18447> A_IWL<18446> A_IWL<18445> A_IWL<18444> A_IWL<18443> A_IWL<18442> A_IWL<18441> A_IWL<18440> A_IWL<18439> A_IWL<18438> A_IWL<18437> A_IWL<18436> A_IWL<18435> A_IWL<18434> A_IWL<18433> A_IWL<18432> A_IWL<19455> A_IWL<19454> A_IWL<19453> A_IWL<19452> A_IWL<19451> A_IWL<19450> A_IWL<19449> A_IWL<19448> A_IWL<19447> A_IWL<19446> A_IWL<19445> A_IWL<19444> A_IWL<19443> A_IWL<19442> A_IWL<19441> A_IWL<19440> A_IWL<19439> A_IWL<19438> A_IWL<19437> A_IWL<19436> A_IWL<19435> A_IWL<19434> A_IWL<19433> A_IWL<19432> A_IWL<19431> A_IWL<19430> A_IWL<19429> A_IWL<19428> A_IWL<19427> A_IWL<19426> A_IWL<19425> A_IWL<19424> A_IWL<19423> A_IWL<19422> A_IWL<19421> A_IWL<19420> A_IWL<19419> A_IWL<19418> A_IWL<19417> A_IWL<19416> A_IWL<19415> A_IWL<19414> A_IWL<19413> A_IWL<19412> A_IWL<19411> A_IWL<19410> A_IWL<19409> A_IWL<19408> A_IWL<19407> A_IWL<19406> A_IWL<19405> A_IWL<19404> A_IWL<19403> A_IWL<19402> A_IWL<19401> A_IWL<19400> A_IWL<19399> A_IWL<19398> A_IWL<19397> A_IWL<19396> A_IWL<19395> A_IWL<19394> A_IWL<19393> A_IWL<19392> A_IWL<19391> A_IWL<19390> A_IWL<19389> A_IWL<19388> A_IWL<19387> A_IWL<19386> A_IWL<19385> A_IWL<19384> A_IWL<19383> A_IWL<19382> A_IWL<19381> A_IWL<19380> A_IWL<19379> A_IWL<19378> A_IWL<19377> A_IWL<19376> A_IWL<19375> A_IWL<19374> A_IWL<19373> A_IWL<19372> A_IWL<19371> A_IWL<19370> A_IWL<19369> A_IWL<19368> A_IWL<19367> A_IWL<19366> A_IWL<19365> A_IWL<19364> A_IWL<19363> A_IWL<19362> A_IWL<19361> A_IWL<19360> A_IWL<19359> A_IWL<19358> A_IWL<19357> A_IWL<19356> A_IWL<19355> A_IWL<19354> A_IWL<19353> A_IWL<19352> A_IWL<19351> A_IWL<19350> A_IWL<19349> A_IWL<19348> A_IWL<19347> A_IWL<19346> A_IWL<19345> A_IWL<19344> A_IWL<19343> A_IWL<19342> A_IWL<19341> A_IWL<19340> A_IWL<19339> A_IWL<19338> A_IWL<19337> A_IWL<19336> A_IWL<19335> A_IWL<19334> A_IWL<19333> A_IWL<19332> A_IWL<19331> A_IWL<19330> A_IWL<19329> A_IWL<19328> A_IWL<19327> A_IWL<19326> A_IWL<19325> A_IWL<19324> A_IWL<19323> A_IWL<19322> A_IWL<19321> A_IWL<19320> A_IWL<19319> A_IWL<19318> A_IWL<19317> A_IWL<19316> A_IWL<19315> A_IWL<19314> A_IWL<19313> A_IWL<19312> A_IWL<19311> A_IWL<19310> A_IWL<19309> A_IWL<19308> A_IWL<19307> A_IWL<19306> A_IWL<19305> A_IWL<19304> A_IWL<19303> A_IWL<19302> A_IWL<19301> A_IWL<19300> A_IWL<19299> A_IWL<19298> A_IWL<19297> A_IWL<19296> A_IWL<19295> A_IWL<19294> A_IWL<19293> A_IWL<19292> A_IWL<19291> A_IWL<19290> A_IWL<19289> A_IWL<19288> A_IWL<19287> A_IWL<19286> A_IWL<19285> A_IWL<19284> A_IWL<19283> A_IWL<19282> A_IWL<19281> A_IWL<19280> A_IWL<19279> A_IWL<19278> A_IWL<19277> A_IWL<19276> A_IWL<19275> A_IWL<19274> A_IWL<19273> A_IWL<19272> A_IWL<19271> A_IWL<19270> A_IWL<19269> A_IWL<19268> A_IWL<19267> A_IWL<19266> A_IWL<19265> A_IWL<19264> A_IWL<19263> A_IWL<19262> A_IWL<19261> A_IWL<19260> A_IWL<19259> A_IWL<19258> A_IWL<19257> A_IWL<19256> A_IWL<19255> A_IWL<19254> A_IWL<19253> A_IWL<19252> A_IWL<19251> A_IWL<19250> A_IWL<19249> A_IWL<19248> A_IWL<19247> A_IWL<19246> A_IWL<19245> A_IWL<19244> A_IWL<19243> A_IWL<19242> A_IWL<19241> A_IWL<19240> A_IWL<19239> A_IWL<19238> A_IWL<19237> A_IWL<19236> A_IWL<19235> A_IWL<19234> A_IWL<19233> A_IWL<19232> A_IWL<19231> A_IWL<19230> A_IWL<19229> A_IWL<19228> A_IWL<19227> A_IWL<19226> A_IWL<19225> A_IWL<19224> A_IWL<19223> A_IWL<19222> A_IWL<19221> A_IWL<19220> A_IWL<19219> A_IWL<19218> A_IWL<19217> A_IWL<19216> A_IWL<19215> A_IWL<19214> A_IWL<19213> A_IWL<19212> A_IWL<19211> A_IWL<19210> A_IWL<19209> A_IWL<19208> A_IWL<19207> A_IWL<19206> A_IWL<19205> A_IWL<19204> A_IWL<19203> A_IWL<19202> A_IWL<19201> A_IWL<19200> A_IWL<19199> A_IWL<19198> A_IWL<19197> A_IWL<19196> A_IWL<19195> A_IWL<19194> A_IWL<19193> A_IWL<19192> A_IWL<19191> A_IWL<19190> A_IWL<19189> A_IWL<19188> A_IWL<19187> A_IWL<19186> A_IWL<19185> A_IWL<19184> A_IWL<19183> A_IWL<19182> A_IWL<19181> A_IWL<19180> A_IWL<19179> A_IWL<19178> A_IWL<19177> A_IWL<19176> A_IWL<19175> A_IWL<19174> A_IWL<19173> A_IWL<19172> A_IWL<19171> A_IWL<19170> A_IWL<19169> A_IWL<19168> A_IWL<19167> A_IWL<19166> A_IWL<19165> A_IWL<19164> A_IWL<19163> A_IWL<19162> A_IWL<19161> A_IWL<19160> A_IWL<19159> A_IWL<19158> A_IWL<19157> A_IWL<19156> A_IWL<19155> A_IWL<19154> A_IWL<19153> A_IWL<19152> A_IWL<19151> A_IWL<19150> A_IWL<19149> A_IWL<19148> A_IWL<19147> A_IWL<19146> A_IWL<19145> A_IWL<19144> A_IWL<19143> A_IWL<19142> A_IWL<19141> A_IWL<19140> A_IWL<19139> A_IWL<19138> A_IWL<19137> A_IWL<19136> A_IWL<19135> A_IWL<19134> A_IWL<19133> A_IWL<19132> A_IWL<19131> A_IWL<19130> A_IWL<19129> A_IWL<19128> A_IWL<19127> A_IWL<19126> A_IWL<19125> A_IWL<19124> A_IWL<19123> A_IWL<19122> A_IWL<19121> A_IWL<19120> A_IWL<19119> A_IWL<19118> A_IWL<19117> A_IWL<19116> A_IWL<19115> A_IWL<19114> A_IWL<19113> A_IWL<19112> A_IWL<19111> A_IWL<19110> A_IWL<19109> A_IWL<19108> A_IWL<19107> A_IWL<19106> A_IWL<19105> A_IWL<19104> A_IWL<19103> A_IWL<19102> A_IWL<19101> A_IWL<19100> A_IWL<19099> A_IWL<19098> A_IWL<19097> A_IWL<19096> A_IWL<19095> A_IWL<19094> A_IWL<19093> A_IWL<19092> A_IWL<19091> A_IWL<19090> A_IWL<19089> A_IWL<19088> A_IWL<19087> A_IWL<19086> A_IWL<19085> A_IWL<19084> A_IWL<19083> A_IWL<19082> A_IWL<19081> A_IWL<19080> A_IWL<19079> A_IWL<19078> A_IWL<19077> A_IWL<19076> A_IWL<19075> A_IWL<19074> A_IWL<19073> A_IWL<19072> A_IWL<19071> A_IWL<19070> A_IWL<19069> A_IWL<19068> A_IWL<19067> A_IWL<19066> A_IWL<19065> A_IWL<19064> A_IWL<19063> A_IWL<19062> A_IWL<19061> A_IWL<19060> A_IWL<19059> A_IWL<19058> A_IWL<19057> A_IWL<19056> A_IWL<19055> A_IWL<19054> A_IWL<19053> A_IWL<19052> A_IWL<19051> A_IWL<19050> A_IWL<19049> A_IWL<19048> A_IWL<19047> A_IWL<19046> A_IWL<19045> A_IWL<19044> A_IWL<19043> A_IWL<19042> A_IWL<19041> A_IWL<19040> A_IWL<19039> A_IWL<19038> A_IWL<19037> A_IWL<19036> A_IWL<19035> A_IWL<19034> A_IWL<19033> A_IWL<19032> A_IWL<19031> A_IWL<19030> A_IWL<19029> A_IWL<19028> A_IWL<19027> A_IWL<19026> A_IWL<19025> A_IWL<19024> A_IWL<19023> A_IWL<19022> A_IWL<19021> A_IWL<19020> A_IWL<19019> A_IWL<19018> A_IWL<19017> A_IWL<19016> A_IWL<19015> A_IWL<19014> A_IWL<19013> A_IWL<19012> A_IWL<19011> A_IWL<19010> A_IWL<19009> A_IWL<19008> A_IWL<19007> A_IWL<19006> A_IWL<19005> A_IWL<19004> A_IWL<19003> A_IWL<19002> A_IWL<19001> A_IWL<19000> A_IWL<18999> A_IWL<18998> A_IWL<18997> A_IWL<18996> A_IWL<18995> A_IWL<18994> A_IWL<18993> A_IWL<18992> A_IWL<18991> A_IWL<18990> A_IWL<18989> A_IWL<18988> A_IWL<18987> A_IWL<18986> A_IWL<18985> A_IWL<18984> A_IWL<18983> A_IWL<18982> A_IWL<18981> A_IWL<18980> A_IWL<18979> A_IWL<18978> A_IWL<18977> A_IWL<18976> A_IWL<18975> A_IWL<18974> A_IWL<18973> A_IWL<18972> A_IWL<18971> A_IWL<18970> A_IWL<18969> A_IWL<18968> A_IWL<18967> A_IWL<18966> A_IWL<18965> A_IWL<18964> A_IWL<18963> A_IWL<18962> A_IWL<18961> A_IWL<18960> A_IWL<18959> A_IWL<18958> A_IWL<18957> A_IWL<18956> A_IWL<18955> A_IWL<18954> A_IWL<18953> A_IWL<18952> A_IWL<18951> A_IWL<18950> A_IWL<18949> A_IWL<18948> A_IWL<18947> A_IWL<18946> A_IWL<18945> A_IWL<18944> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<36> A_BLC<73> A_BLC<72> A_BLC_TOP<73> A_BLC_TOP<72> A_BLT<73> A_BLT<72> A_BLT_TOP<73> A_BLT_TOP<72> A_IWL<18431> A_IWL<18430> A_IWL<18429> A_IWL<18428> A_IWL<18427> A_IWL<18426> A_IWL<18425> A_IWL<18424> A_IWL<18423> A_IWL<18422> A_IWL<18421> A_IWL<18420> A_IWL<18419> A_IWL<18418> A_IWL<18417> A_IWL<18416> A_IWL<18415> A_IWL<18414> A_IWL<18413> A_IWL<18412> A_IWL<18411> A_IWL<18410> A_IWL<18409> A_IWL<18408> A_IWL<18407> A_IWL<18406> A_IWL<18405> A_IWL<18404> A_IWL<18403> A_IWL<18402> A_IWL<18401> A_IWL<18400> A_IWL<18399> A_IWL<18398> A_IWL<18397> A_IWL<18396> A_IWL<18395> A_IWL<18394> A_IWL<18393> A_IWL<18392> A_IWL<18391> A_IWL<18390> A_IWL<18389> A_IWL<18388> A_IWL<18387> A_IWL<18386> A_IWL<18385> A_IWL<18384> A_IWL<18383> A_IWL<18382> A_IWL<18381> A_IWL<18380> A_IWL<18379> A_IWL<18378> A_IWL<18377> A_IWL<18376> A_IWL<18375> A_IWL<18374> A_IWL<18373> A_IWL<18372> A_IWL<18371> A_IWL<18370> A_IWL<18369> A_IWL<18368> A_IWL<18367> A_IWL<18366> A_IWL<18365> A_IWL<18364> A_IWL<18363> A_IWL<18362> A_IWL<18361> A_IWL<18360> A_IWL<18359> A_IWL<18358> A_IWL<18357> A_IWL<18356> A_IWL<18355> A_IWL<18354> A_IWL<18353> A_IWL<18352> A_IWL<18351> A_IWL<18350> A_IWL<18349> A_IWL<18348> A_IWL<18347> A_IWL<18346> A_IWL<18345> A_IWL<18344> A_IWL<18343> A_IWL<18342> A_IWL<18341> A_IWL<18340> A_IWL<18339> A_IWL<18338> A_IWL<18337> A_IWL<18336> A_IWL<18335> A_IWL<18334> A_IWL<18333> A_IWL<18332> A_IWL<18331> A_IWL<18330> A_IWL<18329> A_IWL<18328> A_IWL<18327> A_IWL<18326> A_IWL<18325> A_IWL<18324> A_IWL<18323> A_IWL<18322> A_IWL<18321> A_IWL<18320> A_IWL<18319> A_IWL<18318> A_IWL<18317> A_IWL<18316> A_IWL<18315> A_IWL<18314> A_IWL<18313> A_IWL<18312> A_IWL<18311> A_IWL<18310> A_IWL<18309> A_IWL<18308> A_IWL<18307> A_IWL<18306> A_IWL<18305> A_IWL<18304> A_IWL<18303> A_IWL<18302> A_IWL<18301> A_IWL<18300> A_IWL<18299> A_IWL<18298> A_IWL<18297> A_IWL<18296> A_IWL<18295> A_IWL<18294> A_IWL<18293> A_IWL<18292> A_IWL<18291> A_IWL<18290> A_IWL<18289> A_IWL<18288> A_IWL<18287> A_IWL<18286> A_IWL<18285> A_IWL<18284> A_IWL<18283> A_IWL<18282> A_IWL<18281> A_IWL<18280> A_IWL<18279> A_IWL<18278> A_IWL<18277> A_IWL<18276> A_IWL<18275> A_IWL<18274> A_IWL<18273> A_IWL<18272> A_IWL<18271> A_IWL<18270> A_IWL<18269> A_IWL<18268> A_IWL<18267> A_IWL<18266> A_IWL<18265> A_IWL<18264> A_IWL<18263> A_IWL<18262> A_IWL<18261> A_IWL<18260> A_IWL<18259> A_IWL<18258> A_IWL<18257> A_IWL<18256> A_IWL<18255> A_IWL<18254> A_IWL<18253> A_IWL<18252> A_IWL<18251> A_IWL<18250> A_IWL<18249> A_IWL<18248> A_IWL<18247> A_IWL<18246> A_IWL<18245> A_IWL<18244> A_IWL<18243> A_IWL<18242> A_IWL<18241> A_IWL<18240> A_IWL<18239> A_IWL<18238> A_IWL<18237> A_IWL<18236> A_IWL<18235> A_IWL<18234> A_IWL<18233> A_IWL<18232> A_IWL<18231> A_IWL<18230> A_IWL<18229> A_IWL<18228> A_IWL<18227> A_IWL<18226> A_IWL<18225> A_IWL<18224> A_IWL<18223> A_IWL<18222> A_IWL<18221> A_IWL<18220> A_IWL<18219> A_IWL<18218> A_IWL<18217> A_IWL<18216> A_IWL<18215> A_IWL<18214> A_IWL<18213> A_IWL<18212> A_IWL<18211> A_IWL<18210> A_IWL<18209> A_IWL<18208> A_IWL<18207> A_IWL<18206> A_IWL<18205> A_IWL<18204> A_IWL<18203> A_IWL<18202> A_IWL<18201> A_IWL<18200> A_IWL<18199> A_IWL<18198> A_IWL<18197> A_IWL<18196> A_IWL<18195> A_IWL<18194> A_IWL<18193> A_IWL<18192> A_IWL<18191> A_IWL<18190> A_IWL<18189> A_IWL<18188> A_IWL<18187> A_IWL<18186> A_IWL<18185> A_IWL<18184> A_IWL<18183> A_IWL<18182> A_IWL<18181> A_IWL<18180> A_IWL<18179> A_IWL<18178> A_IWL<18177> A_IWL<18176> A_IWL<18175> A_IWL<18174> A_IWL<18173> A_IWL<18172> A_IWL<18171> A_IWL<18170> A_IWL<18169> A_IWL<18168> A_IWL<18167> A_IWL<18166> A_IWL<18165> A_IWL<18164> A_IWL<18163> A_IWL<18162> A_IWL<18161> A_IWL<18160> A_IWL<18159> A_IWL<18158> A_IWL<18157> A_IWL<18156> A_IWL<18155> A_IWL<18154> A_IWL<18153> A_IWL<18152> A_IWL<18151> A_IWL<18150> A_IWL<18149> A_IWL<18148> A_IWL<18147> A_IWL<18146> A_IWL<18145> A_IWL<18144> A_IWL<18143> A_IWL<18142> A_IWL<18141> A_IWL<18140> A_IWL<18139> A_IWL<18138> A_IWL<18137> A_IWL<18136> A_IWL<18135> A_IWL<18134> A_IWL<18133> A_IWL<18132> A_IWL<18131> A_IWL<18130> A_IWL<18129> A_IWL<18128> A_IWL<18127> A_IWL<18126> A_IWL<18125> A_IWL<18124> A_IWL<18123> A_IWL<18122> A_IWL<18121> A_IWL<18120> A_IWL<18119> A_IWL<18118> A_IWL<18117> A_IWL<18116> A_IWL<18115> A_IWL<18114> A_IWL<18113> A_IWL<18112> A_IWL<18111> A_IWL<18110> A_IWL<18109> A_IWL<18108> A_IWL<18107> A_IWL<18106> A_IWL<18105> A_IWL<18104> A_IWL<18103> A_IWL<18102> A_IWL<18101> A_IWL<18100> A_IWL<18099> A_IWL<18098> A_IWL<18097> A_IWL<18096> A_IWL<18095> A_IWL<18094> A_IWL<18093> A_IWL<18092> A_IWL<18091> A_IWL<18090> A_IWL<18089> A_IWL<18088> A_IWL<18087> A_IWL<18086> A_IWL<18085> A_IWL<18084> A_IWL<18083> A_IWL<18082> A_IWL<18081> A_IWL<18080> A_IWL<18079> A_IWL<18078> A_IWL<18077> A_IWL<18076> A_IWL<18075> A_IWL<18074> A_IWL<18073> A_IWL<18072> A_IWL<18071> A_IWL<18070> A_IWL<18069> A_IWL<18068> A_IWL<18067> A_IWL<18066> A_IWL<18065> A_IWL<18064> A_IWL<18063> A_IWL<18062> A_IWL<18061> A_IWL<18060> A_IWL<18059> A_IWL<18058> A_IWL<18057> A_IWL<18056> A_IWL<18055> A_IWL<18054> A_IWL<18053> A_IWL<18052> A_IWL<18051> A_IWL<18050> A_IWL<18049> A_IWL<18048> A_IWL<18047> A_IWL<18046> A_IWL<18045> A_IWL<18044> A_IWL<18043> A_IWL<18042> A_IWL<18041> A_IWL<18040> A_IWL<18039> A_IWL<18038> A_IWL<18037> A_IWL<18036> A_IWL<18035> A_IWL<18034> A_IWL<18033> A_IWL<18032> A_IWL<18031> A_IWL<18030> A_IWL<18029> A_IWL<18028> A_IWL<18027> A_IWL<18026> A_IWL<18025> A_IWL<18024> A_IWL<18023> A_IWL<18022> A_IWL<18021> A_IWL<18020> A_IWL<18019> A_IWL<18018> A_IWL<18017> A_IWL<18016> A_IWL<18015> A_IWL<18014> A_IWL<18013> A_IWL<18012> A_IWL<18011> A_IWL<18010> A_IWL<18009> A_IWL<18008> A_IWL<18007> A_IWL<18006> A_IWL<18005> A_IWL<18004> A_IWL<18003> A_IWL<18002> A_IWL<18001> A_IWL<18000> A_IWL<17999> A_IWL<17998> A_IWL<17997> A_IWL<17996> A_IWL<17995> A_IWL<17994> A_IWL<17993> A_IWL<17992> A_IWL<17991> A_IWL<17990> A_IWL<17989> A_IWL<17988> A_IWL<17987> A_IWL<17986> A_IWL<17985> A_IWL<17984> A_IWL<17983> A_IWL<17982> A_IWL<17981> A_IWL<17980> A_IWL<17979> A_IWL<17978> A_IWL<17977> A_IWL<17976> A_IWL<17975> A_IWL<17974> A_IWL<17973> A_IWL<17972> A_IWL<17971> A_IWL<17970> A_IWL<17969> A_IWL<17968> A_IWL<17967> A_IWL<17966> A_IWL<17965> A_IWL<17964> A_IWL<17963> A_IWL<17962> A_IWL<17961> A_IWL<17960> A_IWL<17959> A_IWL<17958> A_IWL<17957> A_IWL<17956> A_IWL<17955> A_IWL<17954> A_IWL<17953> A_IWL<17952> A_IWL<17951> A_IWL<17950> A_IWL<17949> A_IWL<17948> A_IWL<17947> A_IWL<17946> A_IWL<17945> A_IWL<17944> A_IWL<17943> A_IWL<17942> A_IWL<17941> A_IWL<17940> A_IWL<17939> A_IWL<17938> A_IWL<17937> A_IWL<17936> A_IWL<17935> A_IWL<17934> A_IWL<17933> A_IWL<17932> A_IWL<17931> A_IWL<17930> A_IWL<17929> A_IWL<17928> A_IWL<17927> A_IWL<17926> A_IWL<17925> A_IWL<17924> A_IWL<17923> A_IWL<17922> A_IWL<17921> A_IWL<17920> A_IWL<18943> A_IWL<18942> A_IWL<18941> A_IWL<18940> A_IWL<18939> A_IWL<18938> A_IWL<18937> A_IWL<18936> A_IWL<18935> A_IWL<18934> A_IWL<18933> A_IWL<18932> A_IWL<18931> A_IWL<18930> A_IWL<18929> A_IWL<18928> A_IWL<18927> A_IWL<18926> A_IWL<18925> A_IWL<18924> A_IWL<18923> A_IWL<18922> A_IWL<18921> A_IWL<18920> A_IWL<18919> A_IWL<18918> A_IWL<18917> A_IWL<18916> A_IWL<18915> A_IWL<18914> A_IWL<18913> A_IWL<18912> A_IWL<18911> A_IWL<18910> A_IWL<18909> A_IWL<18908> A_IWL<18907> A_IWL<18906> A_IWL<18905> A_IWL<18904> A_IWL<18903> A_IWL<18902> A_IWL<18901> A_IWL<18900> A_IWL<18899> A_IWL<18898> A_IWL<18897> A_IWL<18896> A_IWL<18895> A_IWL<18894> A_IWL<18893> A_IWL<18892> A_IWL<18891> A_IWL<18890> A_IWL<18889> A_IWL<18888> A_IWL<18887> A_IWL<18886> A_IWL<18885> A_IWL<18884> A_IWL<18883> A_IWL<18882> A_IWL<18881> A_IWL<18880> A_IWL<18879> A_IWL<18878> A_IWL<18877> A_IWL<18876> A_IWL<18875> A_IWL<18874> A_IWL<18873> A_IWL<18872> A_IWL<18871> A_IWL<18870> A_IWL<18869> A_IWL<18868> A_IWL<18867> A_IWL<18866> A_IWL<18865> A_IWL<18864> A_IWL<18863> A_IWL<18862> A_IWL<18861> A_IWL<18860> A_IWL<18859> A_IWL<18858> A_IWL<18857> A_IWL<18856> A_IWL<18855> A_IWL<18854> A_IWL<18853> A_IWL<18852> A_IWL<18851> A_IWL<18850> A_IWL<18849> A_IWL<18848> A_IWL<18847> A_IWL<18846> A_IWL<18845> A_IWL<18844> A_IWL<18843> A_IWL<18842> A_IWL<18841> A_IWL<18840> A_IWL<18839> A_IWL<18838> A_IWL<18837> A_IWL<18836> A_IWL<18835> A_IWL<18834> A_IWL<18833> A_IWL<18832> A_IWL<18831> A_IWL<18830> A_IWL<18829> A_IWL<18828> A_IWL<18827> A_IWL<18826> A_IWL<18825> A_IWL<18824> A_IWL<18823> A_IWL<18822> A_IWL<18821> A_IWL<18820> A_IWL<18819> A_IWL<18818> A_IWL<18817> A_IWL<18816> A_IWL<18815> A_IWL<18814> A_IWL<18813> A_IWL<18812> A_IWL<18811> A_IWL<18810> A_IWL<18809> A_IWL<18808> A_IWL<18807> A_IWL<18806> A_IWL<18805> A_IWL<18804> A_IWL<18803> A_IWL<18802> A_IWL<18801> A_IWL<18800> A_IWL<18799> A_IWL<18798> A_IWL<18797> A_IWL<18796> A_IWL<18795> A_IWL<18794> A_IWL<18793> A_IWL<18792> A_IWL<18791> A_IWL<18790> A_IWL<18789> A_IWL<18788> A_IWL<18787> A_IWL<18786> A_IWL<18785> A_IWL<18784> A_IWL<18783> A_IWL<18782> A_IWL<18781> A_IWL<18780> A_IWL<18779> A_IWL<18778> A_IWL<18777> A_IWL<18776> A_IWL<18775> A_IWL<18774> A_IWL<18773> A_IWL<18772> A_IWL<18771> A_IWL<18770> A_IWL<18769> A_IWL<18768> A_IWL<18767> A_IWL<18766> A_IWL<18765> A_IWL<18764> A_IWL<18763> A_IWL<18762> A_IWL<18761> A_IWL<18760> A_IWL<18759> A_IWL<18758> A_IWL<18757> A_IWL<18756> A_IWL<18755> A_IWL<18754> A_IWL<18753> A_IWL<18752> A_IWL<18751> A_IWL<18750> A_IWL<18749> A_IWL<18748> A_IWL<18747> A_IWL<18746> A_IWL<18745> A_IWL<18744> A_IWL<18743> A_IWL<18742> A_IWL<18741> A_IWL<18740> A_IWL<18739> A_IWL<18738> A_IWL<18737> A_IWL<18736> A_IWL<18735> A_IWL<18734> A_IWL<18733> A_IWL<18732> A_IWL<18731> A_IWL<18730> A_IWL<18729> A_IWL<18728> A_IWL<18727> A_IWL<18726> A_IWL<18725> A_IWL<18724> A_IWL<18723> A_IWL<18722> A_IWL<18721> A_IWL<18720> A_IWL<18719> A_IWL<18718> A_IWL<18717> A_IWL<18716> A_IWL<18715> A_IWL<18714> A_IWL<18713> A_IWL<18712> A_IWL<18711> A_IWL<18710> A_IWL<18709> A_IWL<18708> A_IWL<18707> A_IWL<18706> A_IWL<18705> A_IWL<18704> A_IWL<18703> A_IWL<18702> A_IWL<18701> A_IWL<18700> A_IWL<18699> A_IWL<18698> A_IWL<18697> A_IWL<18696> A_IWL<18695> A_IWL<18694> A_IWL<18693> A_IWL<18692> A_IWL<18691> A_IWL<18690> A_IWL<18689> A_IWL<18688> A_IWL<18687> A_IWL<18686> A_IWL<18685> A_IWL<18684> A_IWL<18683> A_IWL<18682> A_IWL<18681> A_IWL<18680> A_IWL<18679> A_IWL<18678> A_IWL<18677> A_IWL<18676> A_IWL<18675> A_IWL<18674> A_IWL<18673> A_IWL<18672> A_IWL<18671> A_IWL<18670> A_IWL<18669> A_IWL<18668> A_IWL<18667> A_IWL<18666> A_IWL<18665> A_IWL<18664> A_IWL<18663> A_IWL<18662> A_IWL<18661> A_IWL<18660> A_IWL<18659> A_IWL<18658> A_IWL<18657> A_IWL<18656> A_IWL<18655> A_IWL<18654> A_IWL<18653> A_IWL<18652> A_IWL<18651> A_IWL<18650> A_IWL<18649> A_IWL<18648> A_IWL<18647> A_IWL<18646> A_IWL<18645> A_IWL<18644> A_IWL<18643> A_IWL<18642> A_IWL<18641> A_IWL<18640> A_IWL<18639> A_IWL<18638> A_IWL<18637> A_IWL<18636> A_IWL<18635> A_IWL<18634> A_IWL<18633> A_IWL<18632> A_IWL<18631> A_IWL<18630> A_IWL<18629> A_IWL<18628> A_IWL<18627> A_IWL<18626> A_IWL<18625> A_IWL<18624> A_IWL<18623> A_IWL<18622> A_IWL<18621> A_IWL<18620> A_IWL<18619> A_IWL<18618> A_IWL<18617> A_IWL<18616> A_IWL<18615> A_IWL<18614> A_IWL<18613> A_IWL<18612> A_IWL<18611> A_IWL<18610> A_IWL<18609> A_IWL<18608> A_IWL<18607> A_IWL<18606> A_IWL<18605> A_IWL<18604> A_IWL<18603> A_IWL<18602> A_IWL<18601> A_IWL<18600> A_IWL<18599> A_IWL<18598> A_IWL<18597> A_IWL<18596> A_IWL<18595> A_IWL<18594> A_IWL<18593> A_IWL<18592> A_IWL<18591> A_IWL<18590> A_IWL<18589> A_IWL<18588> A_IWL<18587> A_IWL<18586> A_IWL<18585> A_IWL<18584> A_IWL<18583> A_IWL<18582> A_IWL<18581> A_IWL<18580> A_IWL<18579> A_IWL<18578> A_IWL<18577> A_IWL<18576> A_IWL<18575> A_IWL<18574> A_IWL<18573> A_IWL<18572> A_IWL<18571> A_IWL<18570> A_IWL<18569> A_IWL<18568> A_IWL<18567> A_IWL<18566> A_IWL<18565> A_IWL<18564> A_IWL<18563> A_IWL<18562> A_IWL<18561> A_IWL<18560> A_IWL<18559> A_IWL<18558> A_IWL<18557> A_IWL<18556> A_IWL<18555> A_IWL<18554> A_IWL<18553> A_IWL<18552> A_IWL<18551> A_IWL<18550> A_IWL<18549> A_IWL<18548> A_IWL<18547> A_IWL<18546> A_IWL<18545> A_IWL<18544> A_IWL<18543> A_IWL<18542> A_IWL<18541> A_IWL<18540> A_IWL<18539> A_IWL<18538> A_IWL<18537> A_IWL<18536> A_IWL<18535> A_IWL<18534> A_IWL<18533> A_IWL<18532> A_IWL<18531> A_IWL<18530> A_IWL<18529> A_IWL<18528> A_IWL<18527> A_IWL<18526> A_IWL<18525> A_IWL<18524> A_IWL<18523> A_IWL<18522> A_IWL<18521> A_IWL<18520> A_IWL<18519> A_IWL<18518> A_IWL<18517> A_IWL<18516> A_IWL<18515> A_IWL<18514> A_IWL<18513> A_IWL<18512> A_IWL<18511> A_IWL<18510> A_IWL<18509> A_IWL<18508> A_IWL<18507> A_IWL<18506> A_IWL<18505> A_IWL<18504> A_IWL<18503> A_IWL<18502> A_IWL<18501> A_IWL<18500> A_IWL<18499> A_IWL<18498> A_IWL<18497> A_IWL<18496> A_IWL<18495> A_IWL<18494> A_IWL<18493> A_IWL<18492> A_IWL<18491> A_IWL<18490> A_IWL<18489> A_IWL<18488> A_IWL<18487> A_IWL<18486> A_IWL<18485> A_IWL<18484> A_IWL<18483> A_IWL<18482> A_IWL<18481> A_IWL<18480> A_IWL<18479> A_IWL<18478> A_IWL<18477> A_IWL<18476> A_IWL<18475> A_IWL<18474> A_IWL<18473> A_IWL<18472> A_IWL<18471> A_IWL<18470> A_IWL<18469> A_IWL<18468> A_IWL<18467> A_IWL<18466> A_IWL<18465> A_IWL<18464> A_IWL<18463> A_IWL<18462> A_IWL<18461> A_IWL<18460> A_IWL<18459> A_IWL<18458> A_IWL<18457> A_IWL<18456> A_IWL<18455> A_IWL<18454> A_IWL<18453> A_IWL<18452> A_IWL<18451> A_IWL<18450> A_IWL<18449> A_IWL<18448> A_IWL<18447> A_IWL<18446> A_IWL<18445> A_IWL<18444> A_IWL<18443> A_IWL<18442> A_IWL<18441> A_IWL<18440> A_IWL<18439> A_IWL<18438> A_IWL<18437> A_IWL<18436> A_IWL<18435> A_IWL<18434> A_IWL<18433> A_IWL<18432> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<35> A_BLC<71> A_BLC<70> A_BLC_TOP<71> A_BLC_TOP<70> A_BLT<71> A_BLT<70> A_BLT_TOP<71> A_BLT_TOP<70> A_IWL<17919> A_IWL<17918> A_IWL<17917> A_IWL<17916> A_IWL<17915> A_IWL<17914> A_IWL<17913> A_IWL<17912> A_IWL<17911> A_IWL<17910> A_IWL<17909> A_IWL<17908> A_IWL<17907> A_IWL<17906> A_IWL<17905> A_IWL<17904> A_IWL<17903> A_IWL<17902> A_IWL<17901> A_IWL<17900> A_IWL<17899> A_IWL<17898> A_IWL<17897> A_IWL<17896> A_IWL<17895> A_IWL<17894> A_IWL<17893> A_IWL<17892> A_IWL<17891> A_IWL<17890> A_IWL<17889> A_IWL<17888> A_IWL<17887> A_IWL<17886> A_IWL<17885> A_IWL<17884> A_IWL<17883> A_IWL<17882> A_IWL<17881> A_IWL<17880> A_IWL<17879> A_IWL<17878> A_IWL<17877> A_IWL<17876> A_IWL<17875> A_IWL<17874> A_IWL<17873> A_IWL<17872> A_IWL<17871> A_IWL<17870> A_IWL<17869> A_IWL<17868> A_IWL<17867> A_IWL<17866> A_IWL<17865> A_IWL<17864> A_IWL<17863> A_IWL<17862> A_IWL<17861> A_IWL<17860> A_IWL<17859> A_IWL<17858> A_IWL<17857> A_IWL<17856> A_IWL<17855> A_IWL<17854> A_IWL<17853> A_IWL<17852> A_IWL<17851> A_IWL<17850> A_IWL<17849> A_IWL<17848> A_IWL<17847> A_IWL<17846> A_IWL<17845> A_IWL<17844> A_IWL<17843> A_IWL<17842> A_IWL<17841> A_IWL<17840> A_IWL<17839> A_IWL<17838> A_IWL<17837> A_IWL<17836> A_IWL<17835> A_IWL<17834> A_IWL<17833> A_IWL<17832> A_IWL<17831> A_IWL<17830> A_IWL<17829> A_IWL<17828> A_IWL<17827> A_IWL<17826> A_IWL<17825> A_IWL<17824> A_IWL<17823> A_IWL<17822> A_IWL<17821> A_IWL<17820> A_IWL<17819> A_IWL<17818> A_IWL<17817> A_IWL<17816> A_IWL<17815> A_IWL<17814> A_IWL<17813> A_IWL<17812> A_IWL<17811> A_IWL<17810> A_IWL<17809> A_IWL<17808> A_IWL<17807> A_IWL<17806> A_IWL<17805> A_IWL<17804> A_IWL<17803> A_IWL<17802> A_IWL<17801> A_IWL<17800> A_IWL<17799> A_IWL<17798> A_IWL<17797> A_IWL<17796> A_IWL<17795> A_IWL<17794> A_IWL<17793> A_IWL<17792> A_IWL<17791> A_IWL<17790> A_IWL<17789> A_IWL<17788> A_IWL<17787> A_IWL<17786> A_IWL<17785> A_IWL<17784> A_IWL<17783> A_IWL<17782> A_IWL<17781> A_IWL<17780> A_IWL<17779> A_IWL<17778> A_IWL<17777> A_IWL<17776> A_IWL<17775> A_IWL<17774> A_IWL<17773> A_IWL<17772> A_IWL<17771> A_IWL<17770> A_IWL<17769> A_IWL<17768> A_IWL<17767> A_IWL<17766> A_IWL<17765> A_IWL<17764> A_IWL<17763> A_IWL<17762> A_IWL<17761> A_IWL<17760> A_IWL<17759> A_IWL<17758> A_IWL<17757> A_IWL<17756> A_IWL<17755> A_IWL<17754> A_IWL<17753> A_IWL<17752> A_IWL<17751> A_IWL<17750> A_IWL<17749> A_IWL<17748> A_IWL<17747> A_IWL<17746> A_IWL<17745> A_IWL<17744> A_IWL<17743> A_IWL<17742> A_IWL<17741> A_IWL<17740> A_IWL<17739> A_IWL<17738> A_IWL<17737> A_IWL<17736> A_IWL<17735> A_IWL<17734> A_IWL<17733> A_IWL<17732> A_IWL<17731> A_IWL<17730> A_IWL<17729> A_IWL<17728> A_IWL<17727> A_IWL<17726> A_IWL<17725> A_IWL<17724> A_IWL<17723> A_IWL<17722> A_IWL<17721> A_IWL<17720> A_IWL<17719> A_IWL<17718> A_IWL<17717> A_IWL<17716> A_IWL<17715> A_IWL<17714> A_IWL<17713> A_IWL<17712> A_IWL<17711> A_IWL<17710> A_IWL<17709> A_IWL<17708> A_IWL<17707> A_IWL<17706> A_IWL<17705> A_IWL<17704> A_IWL<17703> A_IWL<17702> A_IWL<17701> A_IWL<17700> A_IWL<17699> A_IWL<17698> A_IWL<17697> A_IWL<17696> A_IWL<17695> A_IWL<17694> A_IWL<17693> A_IWL<17692> A_IWL<17691> A_IWL<17690> A_IWL<17689> A_IWL<17688> A_IWL<17687> A_IWL<17686> A_IWL<17685> A_IWL<17684> A_IWL<17683> A_IWL<17682> A_IWL<17681> A_IWL<17680> A_IWL<17679> A_IWL<17678> A_IWL<17677> A_IWL<17676> A_IWL<17675> A_IWL<17674> A_IWL<17673> A_IWL<17672> A_IWL<17671> A_IWL<17670> A_IWL<17669> A_IWL<17668> A_IWL<17667> A_IWL<17666> A_IWL<17665> A_IWL<17664> A_IWL<17663> A_IWL<17662> A_IWL<17661> A_IWL<17660> A_IWL<17659> A_IWL<17658> A_IWL<17657> A_IWL<17656> A_IWL<17655> A_IWL<17654> A_IWL<17653> A_IWL<17652> A_IWL<17651> A_IWL<17650> A_IWL<17649> A_IWL<17648> A_IWL<17647> A_IWL<17646> A_IWL<17645> A_IWL<17644> A_IWL<17643> A_IWL<17642> A_IWL<17641> A_IWL<17640> A_IWL<17639> A_IWL<17638> A_IWL<17637> A_IWL<17636> A_IWL<17635> A_IWL<17634> A_IWL<17633> A_IWL<17632> A_IWL<17631> A_IWL<17630> A_IWL<17629> A_IWL<17628> A_IWL<17627> A_IWL<17626> A_IWL<17625> A_IWL<17624> A_IWL<17623> A_IWL<17622> A_IWL<17621> A_IWL<17620> A_IWL<17619> A_IWL<17618> A_IWL<17617> A_IWL<17616> A_IWL<17615> A_IWL<17614> A_IWL<17613> A_IWL<17612> A_IWL<17611> A_IWL<17610> A_IWL<17609> A_IWL<17608> A_IWL<17607> A_IWL<17606> A_IWL<17605> A_IWL<17604> A_IWL<17603> A_IWL<17602> A_IWL<17601> A_IWL<17600> A_IWL<17599> A_IWL<17598> A_IWL<17597> A_IWL<17596> A_IWL<17595> A_IWL<17594> A_IWL<17593> A_IWL<17592> A_IWL<17591> A_IWL<17590> A_IWL<17589> A_IWL<17588> A_IWL<17587> A_IWL<17586> A_IWL<17585> A_IWL<17584> A_IWL<17583> A_IWL<17582> A_IWL<17581> A_IWL<17580> A_IWL<17579> A_IWL<17578> A_IWL<17577> A_IWL<17576> A_IWL<17575> A_IWL<17574> A_IWL<17573> A_IWL<17572> A_IWL<17571> A_IWL<17570> A_IWL<17569> A_IWL<17568> A_IWL<17567> A_IWL<17566> A_IWL<17565> A_IWL<17564> A_IWL<17563> A_IWL<17562> A_IWL<17561> A_IWL<17560> A_IWL<17559> A_IWL<17558> A_IWL<17557> A_IWL<17556> A_IWL<17555> A_IWL<17554> A_IWL<17553> A_IWL<17552> A_IWL<17551> A_IWL<17550> A_IWL<17549> A_IWL<17548> A_IWL<17547> A_IWL<17546> A_IWL<17545> A_IWL<17544> A_IWL<17543> A_IWL<17542> A_IWL<17541> A_IWL<17540> A_IWL<17539> A_IWL<17538> A_IWL<17537> A_IWL<17536> A_IWL<17535> A_IWL<17534> A_IWL<17533> A_IWL<17532> A_IWL<17531> A_IWL<17530> A_IWL<17529> A_IWL<17528> A_IWL<17527> A_IWL<17526> A_IWL<17525> A_IWL<17524> A_IWL<17523> A_IWL<17522> A_IWL<17521> A_IWL<17520> A_IWL<17519> A_IWL<17518> A_IWL<17517> A_IWL<17516> A_IWL<17515> A_IWL<17514> A_IWL<17513> A_IWL<17512> A_IWL<17511> A_IWL<17510> A_IWL<17509> A_IWL<17508> A_IWL<17507> A_IWL<17506> A_IWL<17505> A_IWL<17504> A_IWL<17503> A_IWL<17502> A_IWL<17501> A_IWL<17500> A_IWL<17499> A_IWL<17498> A_IWL<17497> A_IWL<17496> A_IWL<17495> A_IWL<17494> A_IWL<17493> A_IWL<17492> A_IWL<17491> A_IWL<17490> A_IWL<17489> A_IWL<17488> A_IWL<17487> A_IWL<17486> A_IWL<17485> A_IWL<17484> A_IWL<17483> A_IWL<17482> A_IWL<17481> A_IWL<17480> A_IWL<17479> A_IWL<17478> A_IWL<17477> A_IWL<17476> A_IWL<17475> A_IWL<17474> A_IWL<17473> A_IWL<17472> A_IWL<17471> A_IWL<17470> A_IWL<17469> A_IWL<17468> A_IWL<17467> A_IWL<17466> A_IWL<17465> A_IWL<17464> A_IWL<17463> A_IWL<17462> A_IWL<17461> A_IWL<17460> A_IWL<17459> A_IWL<17458> A_IWL<17457> A_IWL<17456> A_IWL<17455> A_IWL<17454> A_IWL<17453> A_IWL<17452> A_IWL<17451> A_IWL<17450> A_IWL<17449> A_IWL<17448> A_IWL<17447> A_IWL<17446> A_IWL<17445> A_IWL<17444> A_IWL<17443> A_IWL<17442> A_IWL<17441> A_IWL<17440> A_IWL<17439> A_IWL<17438> A_IWL<17437> A_IWL<17436> A_IWL<17435> A_IWL<17434> A_IWL<17433> A_IWL<17432> A_IWL<17431> A_IWL<17430> A_IWL<17429> A_IWL<17428> A_IWL<17427> A_IWL<17426> A_IWL<17425> A_IWL<17424> A_IWL<17423> A_IWL<17422> A_IWL<17421> A_IWL<17420> A_IWL<17419> A_IWL<17418> A_IWL<17417> A_IWL<17416> A_IWL<17415> A_IWL<17414> A_IWL<17413> A_IWL<17412> A_IWL<17411> A_IWL<17410> A_IWL<17409> A_IWL<17408> A_IWL<18431> A_IWL<18430> A_IWL<18429> A_IWL<18428> A_IWL<18427> A_IWL<18426> A_IWL<18425> A_IWL<18424> A_IWL<18423> A_IWL<18422> A_IWL<18421> A_IWL<18420> A_IWL<18419> A_IWL<18418> A_IWL<18417> A_IWL<18416> A_IWL<18415> A_IWL<18414> A_IWL<18413> A_IWL<18412> A_IWL<18411> A_IWL<18410> A_IWL<18409> A_IWL<18408> A_IWL<18407> A_IWL<18406> A_IWL<18405> A_IWL<18404> A_IWL<18403> A_IWL<18402> A_IWL<18401> A_IWL<18400> A_IWL<18399> A_IWL<18398> A_IWL<18397> A_IWL<18396> A_IWL<18395> A_IWL<18394> A_IWL<18393> A_IWL<18392> A_IWL<18391> A_IWL<18390> A_IWL<18389> A_IWL<18388> A_IWL<18387> A_IWL<18386> A_IWL<18385> A_IWL<18384> A_IWL<18383> A_IWL<18382> A_IWL<18381> A_IWL<18380> A_IWL<18379> A_IWL<18378> A_IWL<18377> A_IWL<18376> A_IWL<18375> A_IWL<18374> A_IWL<18373> A_IWL<18372> A_IWL<18371> A_IWL<18370> A_IWL<18369> A_IWL<18368> A_IWL<18367> A_IWL<18366> A_IWL<18365> A_IWL<18364> A_IWL<18363> A_IWL<18362> A_IWL<18361> A_IWL<18360> A_IWL<18359> A_IWL<18358> A_IWL<18357> A_IWL<18356> A_IWL<18355> A_IWL<18354> A_IWL<18353> A_IWL<18352> A_IWL<18351> A_IWL<18350> A_IWL<18349> A_IWL<18348> A_IWL<18347> A_IWL<18346> A_IWL<18345> A_IWL<18344> A_IWL<18343> A_IWL<18342> A_IWL<18341> A_IWL<18340> A_IWL<18339> A_IWL<18338> A_IWL<18337> A_IWL<18336> A_IWL<18335> A_IWL<18334> A_IWL<18333> A_IWL<18332> A_IWL<18331> A_IWL<18330> A_IWL<18329> A_IWL<18328> A_IWL<18327> A_IWL<18326> A_IWL<18325> A_IWL<18324> A_IWL<18323> A_IWL<18322> A_IWL<18321> A_IWL<18320> A_IWL<18319> A_IWL<18318> A_IWL<18317> A_IWL<18316> A_IWL<18315> A_IWL<18314> A_IWL<18313> A_IWL<18312> A_IWL<18311> A_IWL<18310> A_IWL<18309> A_IWL<18308> A_IWL<18307> A_IWL<18306> A_IWL<18305> A_IWL<18304> A_IWL<18303> A_IWL<18302> A_IWL<18301> A_IWL<18300> A_IWL<18299> A_IWL<18298> A_IWL<18297> A_IWL<18296> A_IWL<18295> A_IWL<18294> A_IWL<18293> A_IWL<18292> A_IWL<18291> A_IWL<18290> A_IWL<18289> A_IWL<18288> A_IWL<18287> A_IWL<18286> A_IWL<18285> A_IWL<18284> A_IWL<18283> A_IWL<18282> A_IWL<18281> A_IWL<18280> A_IWL<18279> A_IWL<18278> A_IWL<18277> A_IWL<18276> A_IWL<18275> A_IWL<18274> A_IWL<18273> A_IWL<18272> A_IWL<18271> A_IWL<18270> A_IWL<18269> A_IWL<18268> A_IWL<18267> A_IWL<18266> A_IWL<18265> A_IWL<18264> A_IWL<18263> A_IWL<18262> A_IWL<18261> A_IWL<18260> A_IWL<18259> A_IWL<18258> A_IWL<18257> A_IWL<18256> A_IWL<18255> A_IWL<18254> A_IWL<18253> A_IWL<18252> A_IWL<18251> A_IWL<18250> A_IWL<18249> A_IWL<18248> A_IWL<18247> A_IWL<18246> A_IWL<18245> A_IWL<18244> A_IWL<18243> A_IWL<18242> A_IWL<18241> A_IWL<18240> A_IWL<18239> A_IWL<18238> A_IWL<18237> A_IWL<18236> A_IWL<18235> A_IWL<18234> A_IWL<18233> A_IWL<18232> A_IWL<18231> A_IWL<18230> A_IWL<18229> A_IWL<18228> A_IWL<18227> A_IWL<18226> A_IWL<18225> A_IWL<18224> A_IWL<18223> A_IWL<18222> A_IWL<18221> A_IWL<18220> A_IWL<18219> A_IWL<18218> A_IWL<18217> A_IWL<18216> A_IWL<18215> A_IWL<18214> A_IWL<18213> A_IWL<18212> A_IWL<18211> A_IWL<18210> A_IWL<18209> A_IWL<18208> A_IWL<18207> A_IWL<18206> A_IWL<18205> A_IWL<18204> A_IWL<18203> A_IWL<18202> A_IWL<18201> A_IWL<18200> A_IWL<18199> A_IWL<18198> A_IWL<18197> A_IWL<18196> A_IWL<18195> A_IWL<18194> A_IWL<18193> A_IWL<18192> A_IWL<18191> A_IWL<18190> A_IWL<18189> A_IWL<18188> A_IWL<18187> A_IWL<18186> A_IWL<18185> A_IWL<18184> A_IWL<18183> A_IWL<18182> A_IWL<18181> A_IWL<18180> A_IWL<18179> A_IWL<18178> A_IWL<18177> A_IWL<18176> A_IWL<18175> A_IWL<18174> A_IWL<18173> A_IWL<18172> A_IWL<18171> A_IWL<18170> A_IWL<18169> A_IWL<18168> A_IWL<18167> A_IWL<18166> A_IWL<18165> A_IWL<18164> A_IWL<18163> A_IWL<18162> A_IWL<18161> A_IWL<18160> A_IWL<18159> A_IWL<18158> A_IWL<18157> A_IWL<18156> A_IWL<18155> A_IWL<18154> A_IWL<18153> A_IWL<18152> A_IWL<18151> A_IWL<18150> A_IWL<18149> A_IWL<18148> A_IWL<18147> A_IWL<18146> A_IWL<18145> A_IWL<18144> A_IWL<18143> A_IWL<18142> A_IWL<18141> A_IWL<18140> A_IWL<18139> A_IWL<18138> A_IWL<18137> A_IWL<18136> A_IWL<18135> A_IWL<18134> A_IWL<18133> A_IWL<18132> A_IWL<18131> A_IWL<18130> A_IWL<18129> A_IWL<18128> A_IWL<18127> A_IWL<18126> A_IWL<18125> A_IWL<18124> A_IWL<18123> A_IWL<18122> A_IWL<18121> A_IWL<18120> A_IWL<18119> A_IWL<18118> A_IWL<18117> A_IWL<18116> A_IWL<18115> A_IWL<18114> A_IWL<18113> A_IWL<18112> A_IWL<18111> A_IWL<18110> A_IWL<18109> A_IWL<18108> A_IWL<18107> A_IWL<18106> A_IWL<18105> A_IWL<18104> A_IWL<18103> A_IWL<18102> A_IWL<18101> A_IWL<18100> A_IWL<18099> A_IWL<18098> A_IWL<18097> A_IWL<18096> A_IWL<18095> A_IWL<18094> A_IWL<18093> A_IWL<18092> A_IWL<18091> A_IWL<18090> A_IWL<18089> A_IWL<18088> A_IWL<18087> A_IWL<18086> A_IWL<18085> A_IWL<18084> A_IWL<18083> A_IWL<18082> A_IWL<18081> A_IWL<18080> A_IWL<18079> A_IWL<18078> A_IWL<18077> A_IWL<18076> A_IWL<18075> A_IWL<18074> A_IWL<18073> A_IWL<18072> A_IWL<18071> A_IWL<18070> A_IWL<18069> A_IWL<18068> A_IWL<18067> A_IWL<18066> A_IWL<18065> A_IWL<18064> A_IWL<18063> A_IWL<18062> A_IWL<18061> A_IWL<18060> A_IWL<18059> A_IWL<18058> A_IWL<18057> A_IWL<18056> A_IWL<18055> A_IWL<18054> A_IWL<18053> A_IWL<18052> A_IWL<18051> A_IWL<18050> A_IWL<18049> A_IWL<18048> A_IWL<18047> A_IWL<18046> A_IWL<18045> A_IWL<18044> A_IWL<18043> A_IWL<18042> A_IWL<18041> A_IWL<18040> A_IWL<18039> A_IWL<18038> A_IWL<18037> A_IWL<18036> A_IWL<18035> A_IWL<18034> A_IWL<18033> A_IWL<18032> A_IWL<18031> A_IWL<18030> A_IWL<18029> A_IWL<18028> A_IWL<18027> A_IWL<18026> A_IWL<18025> A_IWL<18024> A_IWL<18023> A_IWL<18022> A_IWL<18021> A_IWL<18020> A_IWL<18019> A_IWL<18018> A_IWL<18017> A_IWL<18016> A_IWL<18015> A_IWL<18014> A_IWL<18013> A_IWL<18012> A_IWL<18011> A_IWL<18010> A_IWL<18009> A_IWL<18008> A_IWL<18007> A_IWL<18006> A_IWL<18005> A_IWL<18004> A_IWL<18003> A_IWL<18002> A_IWL<18001> A_IWL<18000> A_IWL<17999> A_IWL<17998> A_IWL<17997> A_IWL<17996> A_IWL<17995> A_IWL<17994> A_IWL<17993> A_IWL<17992> A_IWL<17991> A_IWL<17990> A_IWL<17989> A_IWL<17988> A_IWL<17987> A_IWL<17986> A_IWL<17985> A_IWL<17984> A_IWL<17983> A_IWL<17982> A_IWL<17981> A_IWL<17980> A_IWL<17979> A_IWL<17978> A_IWL<17977> A_IWL<17976> A_IWL<17975> A_IWL<17974> A_IWL<17973> A_IWL<17972> A_IWL<17971> A_IWL<17970> A_IWL<17969> A_IWL<17968> A_IWL<17967> A_IWL<17966> A_IWL<17965> A_IWL<17964> A_IWL<17963> A_IWL<17962> A_IWL<17961> A_IWL<17960> A_IWL<17959> A_IWL<17958> A_IWL<17957> A_IWL<17956> A_IWL<17955> A_IWL<17954> A_IWL<17953> A_IWL<17952> A_IWL<17951> A_IWL<17950> A_IWL<17949> A_IWL<17948> A_IWL<17947> A_IWL<17946> A_IWL<17945> A_IWL<17944> A_IWL<17943> A_IWL<17942> A_IWL<17941> A_IWL<17940> A_IWL<17939> A_IWL<17938> A_IWL<17937> A_IWL<17936> A_IWL<17935> A_IWL<17934> A_IWL<17933> A_IWL<17932> A_IWL<17931> A_IWL<17930> A_IWL<17929> A_IWL<17928> A_IWL<17927> A_IWL<17926> A_IWL<17925> A_IWL<17924> A_IWL<17923> A_IWL<17922> A_IWL<17921> A_IWL<17920> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<34> A_BLC<69> A_BLC<68> A_BLC_TOP<69> A_BLC_TOP<68> A_BLT<69> A_BLT<68> A_BLT_TOP<69> A_BLT_TOP<68> A_IWL<17407> A_IWL<17406> A_IWL<17405> A_IWL<17404> A_IWL<17403> A_IWL<17402> A_IWL<17401> A_IWL<17400> A_IWL<17399> A_IWL<17398> A_IWL<17397> A_IWL<17396> A_IWL<17395> A_IWL<17394> A_IWL<17393> A_IWL<17392> A_IWL<17391> A_IWL<17390> A_IWL<17389> A_IWL<17388> A_IWL<17387> A_IWL<17386> A_IWL<17385> A_IWL<17384> A_IWL<17383> A_IWL<17382> A_IWL<17381> A_IWL<17380> A_IWL<17379> A_IWL<17378> A_IWL<17377> A_IWL<17376> A_IWL<17375> A_IWL<17374> A_IWL<17373> A_IWL<17372> A_IWL<17371> A_IWL<17370> A_IWL<17369> A_IWL<17368> A_IWL<17367> A_IWL<17366> A_IWL<17365> A_IWL<17364> A_IWL<17363> A_IWL<17362> A_IWL<17361> A_IWL<17360> A_IWL<17359> A_IWL<17358> A_IWL<17357> A_IWL<17356> A_IWL<17355> A_IWL<17354> A_IWL<17353> A_IWL<17352> A_IWL<17351> A_IWL<17350> A_IWL<17349> A_IWL<17348> A_IWL<17347> A_IWL<17346> A_IWL<17345> A_IWL<17344> A_IWL<17343> A_IWL<17342> A_IWL<17341> A_IWL<17340> A_IWL<17339> A_IWL<17338> A_IWL<17337> A_IWL<17336> A_IWL<17335> A_IWL<17334> A_IWL<17333> A_IWL<17332> A_IWL<17331> A_IWL<17330> A_IWL<17329> A_IWL<17328> A_IWL<17327> A_IWL<17326> A_IWL<17325> A_IWL<17324> A_IWL<17323> A_IWL<17322> A_IWL<17321> A_IWL<17320> A_IWL<17319> A_IWL<17318> A_IWL<17317> A_IWL<17316> A_IWL<17315> A_IWL<17314> A_IWL<17313> A_IWL<17312> A_IWL<17311> A_IWL<17310> A_IWL<17309> A_IWL<17308> A_IWL<17307> A_IWL<17306> A_IWL<17305> A_IWL<17304> A_IWL<17303> A_IWL<17302> A_IWL<17301> A_IWL<17300> A_IWL<17299> A_IWL<17298> A_IWL<17297> A_IWL<17296> A_IWL<17295> A_IWL<17294> A_IWL<17293> A_IWL<17292> A_IWL<17291> A_IWL<17290> A_IWL<17289> A_IWL<17288> A_IWL<17287> A_IWL<17286> A_IWL<17285> A_IWL<17284> A_IWL<17283> A_IWL<17282> A_IWL<17281> A_IWL<17280> A_IWL<17279> A_IWL<17278> A_IWL<17277> A_IWL<17276> A_IWL<17275> A_IWL<17274> A_IWL<17273> A_IWL<17272> A_IWL<17271> A_IWL<17270> A_IWL<17269> A_IWL<17268> A_IWL<17267> A_IWL<17266> A_IWL<17265> A_IWL<17264> A_IWL<17263> A_IWL<17262> A_IWL<17261> A_IWL<17260> A_IWL<17259> A_IWL<17258> A_IWL<17257> A_IWL<17256> A_IWL<17255> A_IWL<17254> A_IWL<17253> A_IWL<17252> A_IWL<17251> A_IWL<17250> A_IWL<17249> A_IWL<17248> A_IWL<17247> A_IWL<17246> A_IWL<17245> A_IWL<17244> A_IWL<17243> A_IWL<17242> A_IWL<17241> A_IWL<17240> A_IWL<17239> A_IWL<17238> A_IWL<17237> A_IWL<17236> A_IWL<17235> A_IWL<17234> A_IWL<17233> A_IWL<17232> A_IWL<17231> A_IWL<17230> A_IWL<17229> A_IWL<17228> A_IWL<17227> A_IWL<17226> A_IWL<17225> A_IWL<17224> A_IWL<17223> A_IWL<17222> A_IWL<17221> A_IWL<17220> A_IWL<17219> A_IWL<17218> A_IWL<17217> A_IWL<17216> A_IWL<17215> A_IWL<17214> A_IWL<17213> A_IWL<17212> A_IWL<17211> A_IWL<17210> A_IWL<17209> A_IWL<17208> A_IWL<17207> A_IWL<17206> A_IWL<17205> A_IWL<17204> A_IWL<17203> A_IWL<17202> A_IWL<17201> A_IWL<17200> A_IWL<17199> A_IWL<17198> A_IWL<17197> A_IWL<17196> A_IWL<17195> A_IWL<17194> A_IWL<17193> A_IWL<17192> A_IWL<17191> A_IWL<17190> A_IWL<17189> A_IWL<17188> A_IWL<17187> A_IWL<17186> A_IWL<17185> A_IWL<17184> A_IWL<17183> A_IWL<17182> A_IWL<17181> A_IWL<17180> A_IWL<17179> A_IWL<17178> A_IWL<17177> A_IWL<17176> A_IWL<17175> A_IWL<17174> A_IWL<17173> A_IWL<17172> A_IWL<17171> A_IWL<17170> A_IWL<17169> A_IWL<17168> A_IWL<17167> A_IWL<17166> A_IWL<17165> A_IWL<17164> A_IWL<17163> A_IWL<17162> A_IWL<17161> A_IWL<17160> A_IWL<17159> A_IWL<17158> A_IWL<17157> A_IWL<17156> A_IWL<17155> A_IWL<17154> A_IWL<17153> A_IWL<17152> A_IWL<17151> A_IWL<17150> A_IWL<17149> A_IWL<17148> A_IWL<17147> A_IWL<17146> A_IWL<17145> A_IWL<17144> A_IWL<17143> A_IWL<17142> A_IWL<17141> A_IWL<17140> A_IWL<17139> A_IWL<17138> A_IWL<17137> A_IWL<17136> A_IWL<17135> A_IWL<17134> A_IWL<17133> A_IWL<17132> A_IWL<17131> A_IWL<17130> A_IWL<17129> A_IWL<17128> A_IWL<17127> A_IWL<17126> A_IWL<17125> A_IWL<17124> A_IWL<17123> A_IWL<17122> A_IWL<17121> A_IWL<17120> A_IWL<17119> A_IWL<17118> A_IWL<17117> A_IWL<17116> A_IWL<17115> A_IWL<17114> A_IWL<17113> A_IWL<17112> A_IWL<17111> A_IWL<17110> A_IWL<17109> A_IWL<17108> A_IWL<17107> A_IWL<17106> A_IWL<17105> A_IWL<17104> A_IWL<17103> A_IWL<17102> A_IWL<17101> A_IWL<17100> A_IWL<17099> A_IWL<17098> A_IWL<17097> A_IWL<17096> A_IWL<17095> A_IWL<17094> A_IWL<17093> A_IWL<17092> A_IWL<17091> A_IWL<17090> A_IWL<17089> A_IWL<17088> A_IWL<17087> A_IWL<17086> A_IWL<17085> A_IWL<17084> A_IWL<17083> A_IWL<17082> A_IWL<17081> A_IWL<17080> A_IWL<17079> A_IWL<17078> A_IWL<17077> A_IWL<17076> A_IWL<17075> A_IWL<17074> A_IWL<17073> A_IWL<17072> A_IWL<17071> A_IWL<17070> A_IWL<17069> A_IWL<17068> A_IWL<17067> A_IWL<17066> A_IWL<17065> A_IWL<17064> A_IWL<17063> A_IWL<17062> A_IWL<17061> A_IWL<17060> A_IWL<17059> A_IWL<17058> A_IWL<17057> A_IWL<17056> A_IWL<17055> A_IWL<17054> A_IWL<17053> A_IWL<17052> A_IWL<17051> A_IWL<17050> A_IWL<17049> A_IWL<17048> A_IWL<17047> A_IWL<17046> A_IWL<17045> A_IWL<17044> A_IWL<17043> A_IWL<17042> A_IWL<17041> A_IWL<17040> A_IWL<17039> A_IWL<17038> A_IWL<17037> A_IWL<17036> A_IWL<17035> A_IWL<17034> A_IWL<17033> A_IWL<17032> A_IWL<17031> A_IWL<17030> A_IWL<17029> A_IWL<17028> A_IWL<17027> A_IWL<17026> A_IWL<17025> A_IWL<17024> A_IWL<17023> A_IWL<17022> A_IWL<17021> A_IWL<17020> A_IWL<17019> A_IWL<17018> A_IWL<17017> A_IWL<17016> A_IWL<17015> A_IWL<17014> A_IWL<17013> A_IWL<17012> A_IWL<17011> A_IWL<17010> A_IWL<17009> A_IWL<17008> A_IWL<17007> A_IWL<17006> A_IWL<17005> A_IWL<17004> A_IWL<17003> A_IWL<17002> A_IWL<17001> A_IWL<17000> A_IWL<16999> A_IWL<16998> A_IWL<16997> A_IWL<16996> A_IWL<16995> A_IWL<16994> A_IWL<16993> A_IWL<16992> A_IWL<16991> A_IWL<16990> A_IWL<16989> A_IWL<16988> A_IWL<16987> A_IWL<16986> A_IWL<16985> A_IWL<16984> A_IWL<16983> A_IWL<16982> A_IWL<16981> A_IWL<16980> A_IWL<16979> A_IWL<16978> A_IWL<16977> A_IWL<16976> A_IWL<16975> A_IWL<16974> A_IWL<16973> A_IWL<16972> A_IWL<16971> A_IWL<16970> A_IWL<16969> A_IWL<16968> A_IWL<16967> A_IWL<16966> A_IWL<16965> A_IWL<16964> A_IWL<16963> A_IWL<16962> A_IWL<16961> A_IWL<16960> A_IWL<16959> A_IWL<16958> A_IWL<16957> A_IWL<16956> A_IWL<16955> A_IWL<16954> A_IWL<16953> A_IWL<16952> A_IWL<16951> A_IWL<16950> A_IWL<16949> A_IWL<16948> A_IWL<16947> A_IWL<16946> A_IWL<16945> A_IWL<16944> A_IWL<16943> A_IWL<16942> A_IWL<16941> A_IWL<16940> A_IWL<16939> A_IWL<16938> A_IWL<16937> A_IWL<16936> A_IWL<16935> A_IWL<16934> A_IWL<16933> A_IWL<16932> A_IWL<16931> A_IWL<16930> A_IWL<16929> A_IWL<16928> A_IWL<16927> A_IWL<16926> A_IWL<16925> A_IWL<16924> A_IWL<16923> A_IWL<16922> A_IWL<16921> A_IWL<16920> A_IWL<16919> A_IWL<16918> A_IWL<16917> A_IWL<16916> A_IWL<16915> A_IWL<16914> A_IWL<16913> A_IWL<16912> A_IWL<16911> A_IWL<16910> A_IWL<16909> A_IWL<16908> A_IWL<16907> A_IWL<16906> A_IWL<16905> A_IWL<16904> A_IWL<16903> A_IWL<16902> A_IWL<16901> A_IWL<16900> A_IWL<16899> A_IWL<16898> A_IWL<16897> A_IWL<16896> A_IWL<17919> A_IWL<17918> A_IWL<17917> A_IWL<17916> A_IWL<17915> A_IWL<17914> A_IWL<17913> A_IWL<17912> A_IWL<17911> A_IWL<17910> A_IWL<17909> A_IWL<17908> A_IWL<17907> A_IWL<17906> A_IWL<17905> A_IWL<17904> A_IWL<17903> A_IWL<17902> A_IWL<17901> A_IWL<17900> A_IWL<17899> A_IWL<17898> A_IWL<17897> A_IWL<17896> A_IWL<17895> A_IWL<17894> A_IWL<17893> A_IWL<17892> A_IWL<17891> A_IWL<17890> A_IWL<17889> A_IWL<17888> A_IWL<17887> A_IWL<17886> A_IWL<17885> A_IWL<17884> A_IWL<17883> A_IWL<17882> A_IWL<17881> A_IWL<17880> A_IWL<17879> A_IWL<17878> A_IWL<17877> A_IWL<17876> A_IWL<17875> A_IWL<17874> A_IWL<17873> A_IWL<17872> A_IWL<17871> A_IWL<17870> A_IWL<17869> A_IWL<17868> A_IWL<17867> A_IWL<17866> A_IWL<17865> A_IWL<17864> A_IWL<17863> A_IWL<17862> A_IWL<17861> A_IWL<17860> A_IWL<17859> A_IWL<17858> A_IWL<17857> A_IWL<17856> A_IWL<17855> A_IWL<17854> A_IWL<17853> A_IWL<17852> A_IWL<17851> A_IWL<17850> A_IWL<17849> A_IWL<17848> A_IWL<17847> A_IWL<17846> A_IWL<17845> A_IWL<17844> A_IWL<17843> A_IWL<17842> A_IWL<17841> A_IWL<17840> A_IWL<17839> A_IWL<17838> A_IWL<17837> A_IWL<17836> A_IWL<17835> A_IWL<17834> A_IWL<17833> A_IWL<17832> A_IWL<17831> A_IWL<17830> A_IWL<17829> A_IWL<17828> A_IWL<17827> A_IWL<17826> A_IWL<17825> A_IWL<17824> A_IWL<17823> A_IWL<17822> A_IWL<17821> A_IWL<17820> A_IWL<17819> A_IWL<17818> A_IWL<17817> A_IWL<17816> A_IWL<17815> A_IWL<17814> A_IWL<17813> A_IWL<17812> A_IWL<17811> A_IWL<17810> A_IWL<17809> A_IWL<17808> A_IWL<17807> A_IWL<17806> A_IWL<17805> A_IWL<17804> A_IWL<17803> A_IWL<17802> A_IWL<17801> A_IWL<17800> A_IWL<17799> A_IWL<17798> A_IWL<17797> A_IWL<17796> A_IWL<17795> A_IWL<17794> A_IWL<17793> A_IWL<17792> A_IWL<17791> A_IWL<17790> A_IWL<17789> A_IWL<17788> A_IWL<17787> A_IWL<17786> A_IWL<17785> A_IWL<17784> A_IWL<17783> A_IWL<17782> A_IWL<17781> A_IWL<17780> A_IWL<17779> A_IWL<17778> A_IWL<17777> A_IWL<17776> A_IWL<17775> A_IWL<17774> A_IWL<17773> A_IWL<17772> A_IWL<17771> A_IWL<17770> A_IWL<17769> A_IWL<17768> A_IWL<17767> A_IWL<17766> A_IWL<17765> A_IWL<17764> A_IWL<17763> A_IWL<17762> A_IWL<17761> A_IWL<17760> A_IWL<17759> A_IWL<17758> A_IWL<17757> A_IWL<17756> A_IWL<17755> A_IWL<17754> A_IWL<17753> A_IWL<17752> A_IWL<17751> A_IWL<17750> A_IWL<17749> A_IWL<17748> A_IWL<17747> A_IWL<17746> A_IWL<17745> A_IWL<17744> A_IWL<17743> A_IWL<17742> A_IWL<17741> A_IWL<17740> A_IWL<17739> A_IWL<17738> A_IWL<17737> A_IWL<17736> A_IWL<17735> A_IWL<17734> A_IWL<17733> A_IWL<17732> A_IWL<17731> A_IWL<17730> A_IWL<17729> A_IWL<17728> A_IWL<17727> A_IWL<17726> A_IWL<17725> A_IWL<17724> A_IWL<17723> A_IWL<17722> A_IWL<17721> A_IWL<17720> A_IWL<17719> A_IWL<17718> A_IWL<17717> A_IWL<17716> A_IWL<17715> A_IWL<17714> A_IWL<17713> A_IWL<17712> A_IWL<17711> A_IWL<17710> A_IWL<17709> A_IWL<17708> A_IWL<17707> A_IWL<17706> A_IWL<17705> A_IWL<17704> A_IWL<17703> A_IWL<17702> A_IWL<17701> A_IWL<17700> A_IWL<17699> A_IWL<17698> A_IWL<17697> A_IWL<17696> A_IWL<17695> A_IWL<17694> A_IWL<17693> A_IWL<17692> A_IWL<17691> A_IWL<17690> A_IWL<17689> A_IWL<17688> A_IWL<17687> A_IWL<17686> A_IWL<17685> A_IWL<17684> A_IWL<17683> A_IWL<17682> A_IWL<17681> A_IWL<17680> A_IWL<17679> A_IWL<17678> A_IWL<17677> A_IWL<17676> A_IWL<17675> A_IWL<17674> A_IWL<17673> A_IWL<17672> A_IWL<17671> A_IWL<17670> A_IWL<17669> A_IWL<17668> A_IWL<17667> A_IWL<17666> A_IWL<17665> A_IWL<17664> A_IWL<17663> A_IWL<17662> A_IWL<17661> A_IWL<17660> A_IWL<17659> A_IWL<17658> A_IWL<17657> A_IWL<17656> A_IWL<17655> A_IWL<17654> A_IWL<17653> A_IWL<17652> A_IWL<17651> A_IWL<17650> A_IWL<17649> A_IWL<17648> A_IWL<17647> A_IWL<17646> A_IWL<17645> A_IWL<17644> A_IWL<17643> A_IWL<17642> A_IWL<17641> A_IWL<17640> A_IWL<17639> A_IWL<17638> A_IWL<17637> A_IWL<17636> A_IWL<17635> A_IWL<17634> A_IWL<17633> A_IWL<17632> A_IWL<17631> A_IWL<17630> A_IWL<17629> A_IWL<17628> A_IWL<17627> A_IWL<17626> A_IWL<17625> A_IWL<17624> A_IWL<17623> A_IWL<17622> A_IWL<17621> A_IWL<17620> A_IWL<17619> A_IWL<17618> A_IWL<17617> A_IWL<17616> A_IWL<17615> A_IWL<17614> A_IWL<17613> A_IWL<17612> A_IWL<17611> A_IWL<17610> A_IWL<17609> A_IWL<17608> A_IWL<17607> A_IWL<17606> A_IWL<17605> A_IWL<17604> A_IWL<17603> A_IWL<17602> A_IWL<17601> A_IWL<17600> A_IWL<17599> A_IWL<17598> A_IWL<17597> A_IWL<17596> A_IWL<17595> A_IWL<17594> A_IWL<17593> A_IWL<17592> A_IWL<17591> A_IWL<17590> A_IWL<17589> A_IWL<17588> A_IWL<17587> A_IWL<17586> A_IWL<17585> A_IWL<17584> A_IWL<17583> A_IWL<17582> A_IWL<17581> A_IWL<17580> A_IWL<17579> A_IWL<17578> A_IWL<17577> A_IWL<17576> A_IWL<17575> A_IWL<17574> A_IWL<17573> A_IWL<17572> A_IWL<17571> A_IWL<17570> A_IWL<17569> A_IWL<17568> A_IWL<17567> A_IWL<17566> A_IWL<17565> A_IWL<17564> A_IWL<17563> A_IWL<17562> A_IWL<17561> A_IWL<17560> A_IWL<17559> A_IWL<17558> A_IWL<17557> A_IWL<17556> A_IWL<17555> A_IWL<17554> A_IWL<17553> A_IWL<17552> A_IWL<17551> A_IWL<17550> A_IWL<17549> A_IWL<17548> A_IWL<17547> A_IWL<17546> A_IWL<17545> A_IWL<17544> A_IWL<17543> A_IWL<17542> A_IWL<17541> A_IWL<17540> A_IWL<17539> A_IWL<17538> A_IWL<17537> A_IWL<17536> A_IWL<17535> A_IWL<17534> A_IWL<17533> A_IWL<17532> A_IWL<17531> A_IWL<17530> A_IWL<17529> A_IWL<17528> A_IWL<17527> A_IWL<17526> A_IWL<17525> A_IWL<17524> A_IWL<17523> A_IWL<17522> A_IWL<17521> A_IWL<17520> A_IWL<17519> A_IWL<17518> A_IWL<17517> A_IWL<17516> A_IWL<17515> A_IWL<17514> A_IWL<17513> A_IWL<17512> A_IWL<17511> A_IWL<17510> A_IWL<17509> A_IWL<17508> A_IWL<17507> A_IWL<17506> A_IWL<17505> A_IWL<17504> A_IWL<17503> A_IWL<17502> A_IWL<17501> A_IWL<17500> A_IWL<17499> A_IWL<17498> A_IWL<17497> A_IWL<17496> A_IWL<17495> A_IWL<17494> A_IWL<17493> A_IWL<17492> A_IWL<17491> A_IWL<17490> A_IWL<17489> A_IWL<17488> A_IWL<17487> A_IWL<17486> A_IWL<17485> A_IWL<17484> A_IWL<17483> A_IWL<17482> A_IWL<17481> A_IWL<17480> A_IWL<17479> A_IWL<17478> A_IWL<17477> A_IWL<17476> A_IWL<17475> A_IWL<17474> A_IWL<17473> A_IWL<17472> A_IWL<17471> A_IWL<17470> A_IWL<17469> A_IWL<17468> A_IWL<17467> A_IWL<17466> A_IWL<17465> A_IWL<17464> A_IWL<17463> A_IWL<17462> A_IWL<17461> A_IWL<17460> A_IWL<17459> A_IWL<17458> A_IWL<17457> A_IWL<17456> A_IWL<17455> A_IWL<17454> A_IWL<17453> A_IWL<17452> A_IWL<17451> A_IWL<17450> A_IWL<17449> A_IWL<17448> A_IWL<17447> A_IWL<17446> A_IWL<17445> A_IWL<17444> A_IWL<17443> A_IWL<17442> A_IWL<17441> A_IWL<17440> A_IWL<17439> A_IWL<17438> A_IWL<17437> A_IWL<17436> A_IWL<17435> A_IWL<17434> A_IWL<17433> A_IWL<17432> A_IWL<17431> A_IWL<17430> A_IWL<17429> A_IWL<17428> A_IWL<17427> A_IWL<17426> A_IWL<17425> A_IWL<17424> A_IWL<17423> A_IWL<17422> A_IWL<17421> A_IWL<17420> A_IWL<17419> A_IWL<17418> A_IWL<17417> A_IWL<17416> A_IWL<17415> A_IWL<17414> A_IWL<17413> A_IWL<17412> A_IWL<17411> A_IWL<17410> A_IWL<17409> A_IWL<17408> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<33> A_BLC<67> A_BLC<66> A_BLC_TOP<67> A_BLC_TOP<66> A_BLT<67> A_BLT<66> A_BLT_TOP<67> A_BLT_TOP<66> A_IWL<16895> A_IWL<16894> A_IWL<16893> A_IWL<16892> A_IWL<16891> A_IWL<16890> A_IWL<16889> A_IWL<16888> A_IWL<16887> A_IWL<16886> A_IWL<16885> A_IWL<16884> A_IWL<16883> A_IWL<16882> A_IWL<16881> A_IWL<16880> A_IWL<16879> A_IWL<16878> A_IWL<16877> A_IWL<16876> A_IWL<16875> A_IWL<16874> A_IWL<16873> A_IWL<16872> A_IWL<16871> A_IWL<16870> A_IWL<16869> A_IWL<16868> A_IWL<16867> A_IWL<16866> A_IWL<16865> A_IWL<16864> A_IWL<16863> A_IWL<16862> A_IWL<16861> A_IWL<16860> A_IWL<16859> A_IWL<16858> A_IWL<16857> A_IWL<16856> A_IWL<16855> A_IWL<16854> A_IWL<16853> A_IWL<16852> A_IWL<16851> A_IWL<16850> A_IWL<16849> A_IWL<16848> A_IWL<16847> A_IWL<16846> A_IWL<16845> A_IWL<16844> A_IWL<16843> A_IWL<16842> A_IWL<16841> A_IWL<16840> A_IWL<16839> A_IWL<16838> A_IWL<16837> A_IWL<16836> A_IWL<16835> A_IWL<16834> A_IWL<16833> A_IWL<16832> A_IWL<16831> A_IWL<16830> A_IWL<16829> A_IWL<16828> A_IWL<16827> A_IWL<16826> A_IWL<16825> A_IWL<16824> A_IWL<16823> A_IWL<16822> A_IWL<16821> A_IWL<16820> A_IWL<16819> A_IWL<16818> A_IWL<16817> A_IWL<16816> A_IWL<16815> A_IWL<16814> A_IWL<16813> A_IWL<16812> A_IWL<16811> A_IWL<16810> A_IWL<16809> A_IWL<16808> A_IWL<16807> A_IWL<16806> A_IWL<16805> A_IWL<16804> A_IWL<16803> A_IWL<16802> A_IWL<16801> A_IWL<16800> A_IWL<16799> A_IWL<16798> A_IWL<16797> A_IWL<16796> A_IWL<16795> A_IWL<16794> A_IWL<16793> A_IWL<16792> A_IWL<16791> A_IWL<16790> A_IWL<16789> A_IWL<16788> A_IWL<16787> A_IWL<16786> A_IWL<16785> A_IWL<16784> A_IWL<16783> A_IWL<16782> A_IWL<16781> A_IWL<16780> A_IWL<16779> A_IWL<16778> A_IWL<16777> A_IWL<16776> A_IWL<16775> A_IWL<16774> A_IWL<16773> A_IWL<16772> A_IWL<16771> A_IWL<16770> A_IWL<16769> A_IWL<16768> A_IWL<16767> A_IWL<16766> A_IWL<16765> A_IWL<16764> A_IWL<16763> A_IWL<16762> A_IWL<16761> A_IWL<16760> A_IWL<16759> A_IWL<16758> A_IWL<16757> A_IWL<16756> A_IWL<16755> A_IWL<16754> A_IWL<16753> A_IWL<16752> A_IWL<16751> A_IWL<16750> A_IWL<16749> A_IWL<16748> A_IWL<16747> A_IWL<16746> A_IWL<16745> A_IWL<16744> A_IWL<16743> A_IWL<16742> A_IWL<16741> A_IWL<16740> A_IWL<16739> A_IWL<16738> A_IWL<16737> A_IWL<16736> A_IWL<16735> A_IWL<16734> A_IWL<16733> A_IWL<16732> A_IWL<16731> A_IWL<16730> A_IWL<16729> A_IWL<16728> A_IWL<16727> A_IWL<16726> A_IWL<16725> A_IWL<16724> A_IWL<16723> A_IWL<16722> A_IWL<16721> A_IWL<16720> A_IWL<16719> A_IWL<16718> A_IWL<16717> A_IWL<16716> A_IWL<16715> A_IWL<16714> A_IWL<16713> A_IWL<16712> A_IWL<16711> A_IWL<16710> A_IWL<16709> A_IWL<16708> A_IWL<16707> A_IWL<16706> A_IWL<16705> A_IWL<16704> A_IWL<16703> A_IWL<16702> A_IWL<16701> A_IWL<16700> A_IWL<16699> A_IWL<16698> A_IWL<16697> A_IWL<16696> A_IWL<16695> A_IWL<16694> A_IWL<16693> A_IWL<16692> A_IWL<16691> A_IWL<16690> A_IWL<16689> A_IWL<16688> A_IWL<16687> A_IWL<16686> A_IWL<16685> A_IWL<16684> A_IWL<16683> A_IWL<16682> A_IWL<16681> A_IWL<16680> A_IWL<16679> A_IWL<16678> A_IWL<16677> A_IWL<16676> A_IWL<16675> A_IWL<16674> A_IWL<16673> A_IWL<16672> A_IWL<16671> A_IWL<16670> A_IWL<16669> A_IWL<16668> A_IWL<16667> A_IWL<16666> A_IWL<16665> A_IWL<16664> A_IWL<16663> A_IWL<16662> A_IWL<16661> A_IWL<16660> A_IWL<16659> A_IWL<16658> A_IWL<16657> A_IWL<16656> A_IWL<16655> A_IWL<16654> A_IWL<16653> A_IWL<16652> A_IWL<16651> A_IWL<16650> A_IWL<16649> A_IWL<16648> A_IWL<16647> A_IWL<16646> A_IWL<16645> A_IWL<16644> A_IWL<16643> A_IWL<16642> A_IWL<16641> A_IWL<16640> A_IWL<16639> A_IWL<16638> A_IWL<16637> A_IWL<16636> A_IWL<16635> A_IWL<16634> A_IWL<16633> A_IWL<16632> A_IWL<16631> A_IWL<16630> A_IWL<16629> A_IWL<16628> A_IWL<16627> A_IWL<16626> A_IWL<16625> A_IWL<16624> A_IWL<16623> A_IWL<16622> A_IWL<16621> A_IWL<16620> A_IWL<16619> A_IWL<16618> A_IWL<16617> A_IWL<16616> A_IWL<16615> A_IWL<16614> A_IWL<16613> A_IWL<16612> A_IWL<16611> A_IWL<16610> A_IWL<16609> A_IWL<16608> A_IWL<16607> A_IWL<16606> A_IWL<16605> A_IWL<16604> A_IWL<16603> A_IWL<16602> A_IWL<16601> A_IWL<16600> A_IWL<16599> A_IWL<16598> A_IWL<16597> A_IWL<16596> A_IWL<16595> A_IWL<16594> A_IWL<16593> A_IWL<16592> A_IWL<16591> A_IWL<16590> A_IWL<16589> A_IWL<16588> A_IWL<16587> A_IWL<16586> A_IWL<16585> A_IWL<16584> A_IWL<16583> A_IWL<16582> A_IWL<16581> A_IWL<16580> A_IWL<16579> A_IWL<16578> A_IWL<16577> A_IWL<16576> A_IWL<16575> A_IWL<16574> A_IWL<16573> A_IWL<16572> A_IWL<16571> A_IWL<16570> A_IWL<16569> A_IWL<16568> A_IWL<16567> A_IWL<16566> A_IWL<16565> A_IWL<16564> A_IWL<16563> A_IWL<16562> A_IWL<16561> A_IWL<16560> A_IWL<16559> A_IWL<16558> A_IWL<16557> A_IWL<16556> A_IWL<16555> A_IWL<16554> A_IWL<16553> A_IWL<16552> A_IWL<16551> A_IWL<16550> A_IWL<16549> A_IWL<16548> A_IWL<16547> A_IWL<16546> A_IWL<16545> A_IWL<16544> A_IWL<16543> A_IWL<16542> A_IWL<16541> A_IWL<16540> A_IWL<16539> A_IWL<16538> A_IWL<16537> A_IWL<16536> A_IWL<16535> A_IWL<16534> A_IWL<16533> A_IWL<16532> A_IWL<16531> A_IWL<16530> A_IWL<16529> A_IWL<16528> A_IWL<16527> A_IWL<16526> A_IWL<16525> A_IWL<16524> A_IWL<16523> A_IWL<16522> A_IWL<16521> A_IWL<16520> A_IWL<16519> A_IWL<16518> A_IWL<16517> A_IWL<16516> A_IWL<16515> A_IWL<16514> A_IWL<16513> A_IWL<16512> A_IWL<16511> A_IWL<16510> A_IWL<16509> A_IWL<16508> A_IWL<16507> A_IWL<16506> A_IWL<16505> A_IWL<16504> A_IWL<16503> A_IWL<16502> A_IWL<16501> A_IWL<16500> A_IWL<16499> A_IWL<16498> A_IWL<16497> A_IWL<16496> A_IWL<16495> A_IWL<16494> A_IWL<16493> A_IWL<16492> A_IWL<16491> A_IWL<16490> A_IWL<16489> A_IWL<16488> A_IWL<16487> A_IWL<16486> A_IWL<16485> A_IWL<16484> A_IWL<16483> A_IWL<16482> A_IWL<16481> A_IWL<16480> A_IWL<16479> A_IWL<16478> A_IWL<16477> A_IWL<16476> A_IWL<16475> A_IWL<16474> A_IWL<16473> A_IWL<16472> A_IWL<16471> A_IWL<16470> A_IWL<16469> A_IWL<16468> A_IWL<16467> A_IWL<16466> A_IWL<16465> A_IWL<16464> A_IWL<16463> A_IWL<16462> A_IWL<16461> A_IWL<16460> A_IWL<16459> A_IWL<16458> A_IWL<16457> A_IWL<16456> A_IWL<16455> A_IWL<16454> A_IWL<16453> A_IWL<16452> A_IWL<16451> A_IWL<16450> A_IWL<16449> A_IWL<16448> A_IWL<16447> A_IWL<16446> A_IWL<16445> A_IWL<16444> A_IWL<16443> A_IWL<16442> A_IWL<16441> A_IWL<16440> A_IWL<16439> A_IWL<16438> A_IWL<16437> A_IWL<16436> A_IWL<16435> A_IWL<16434> A_IWL<16433> A_IWL<16432> A_IWL<16431> A_IWL<16430> A_IWL<16429> A_IWL<16428> A_IWL<16427> A_IWL<16426> A_IWL<16425> A_IWL<16424> A_IWL<16423> A_IWL<16422> A_IWL<16421> A_IWL<16420> A_IWL<16419> A_IWL<16418> A_IWL<16417> A_IWL<16416> A_IWL<16415> A_IWL<16414> A_IWL<16413> A_IWL<16412> A_IWL<16411> A_IWL<16410> A_IWL<16409> A_IWL<16408> A_IWL<16407> A_IWL<16406> A_IWL<16405> A_IWL<16404> A_IWL<16403> A_IWL<16402> A_IWL<16401> A_IWL<16400> A_IWL<16399> A_IWL<16398> A_IWL<16397> A_IWL<16396> A_IWL<16395> A_IWL<16394> A_IWL<16393> A_IWL<16392> A_IWL<16391> A_IWL<16390> A_IWL<16389> A_IWL<16388> A_IWL<16387> A_IWL<16386> A_IWL<16385> A_IWL<16384> A_IWL<17407> A_IWL<17406> A_IWL<17405> A_IWL<17404> A_IWL<17403> A_IWL<17402> A_IWL<17401> A_IWL<17400> A_IWL<17399> A_IWL<17398> A_IWL<17397> A_IWL<17396> A_IWL<17395> A_IWL<17394> A_IWL<17393> A_IWL<17392> A_IWL<17391> A_IWL<17390> A_IWL<17389> A_IWL<17388> A_IWL<17387> A_IWL<17386> A_IWL<17385> A_IWL<17384> A_IWL<17383> A_IWL<17382> A_IWL<17381> A_IWL<17380> A_IWL<17379> A_IWL<17378> A_IWL<17377> A_IWL<17376> A_IWL<17375> A_IWL<17374> A_IWL<17373> A_IWL<17372> A_IWL<17371> A_IWL<17370> A_IWL<17369> A_IWL<17368> A_IWL<17367> A_IWL<17366> A_IWL<17365> A_IWL<17364> A_IWL<17363> A_IWL<17362> A_IWL<17361> A_IWL<17360> A_IWL<17359> A_IWL<17358> A_IWL<17357> A_IWL<17356> A_IWL<17355> A_IWL<17354> A_IWL<17353> A_IWL<17352> A_IWL<17351> A_IWL<17350> A_IWL<17349> A_IWL<17348> A_IWL<17347> A_IWL<17346> A_IWL<17345> A_IWL<17344> A_IWL<17343> A_IWL<17342> A_IWL<17341> A_IWL<17340> A_IWL<17339> A_IWL<17338> A_IWL<17337> A_IWL<17336> A_IWL<17335> A_IWL<17334> A_IWL<17333> A_IWL<17332> A_IWL<17331> A_IWL<17330> A_IWL<17329> A_IWL<17328> A_IWL<17327> A_IWL<17326> A_IWL<17325> A_IWL<17324> A_IWL<17323> A_IWL<17322> A_IWL<17321> A_IWL<17320> A_IWL<17319> A_IWL<17318> A_IWL<17317> A_IWL<17316> A_IWL<17315> A_IWL<17314> A_IWL<17313> A_IWL<17312> A_IWL<17311> A_IWL<17310> A_IWL<17309> A_IWL<17308> A_IWL<17307> A_IWL<17306> A_IWL<17305> A_IWL<17304> A_IWL<17303> A_IWL<17302> A_IWL<17301> A_IWL<17300> A_IWL<17299> A_IWL<17298> A_IWL<17297> A_IWL<17296> A_IWL<17295> A_IWL<17294> A_IWL<17293> A_IWL<17292> A_IWL<17291> A_IWL<17290> A_IWL<17289> A_IWL<17288> A_IWL<17287> A_IWL<17286> A_IWL<17285> A_IWL<17284> A_IWL<17283> A_IWL<17282> A_IWL<17281> A_IWL<17280> A_IWL<17279> A_IWL<17278> A_IWL<17277> A_IWL<17276> A_IWL<17275> A_IWL<17274> A_IWL<17273> A_IWL<17272> A_IWL<17271> A_IWL<17270> A_IWL<17269> A_IWL<17268> A_IWL<17267> A_IWL<17266> A_IWL<17265> A_IWL<17264> A_IWL<17263> A_IWL<17262> A_IWL<17261> A_IWL<17260> A_IWL<17259> A_IWL<17258> A_IWL<17257> A_IWL<17256> A_IWL<17255> A_IWL<17254> A_IWL<17253> A_IWL<17252> A_IWL<17251> A_IWL<17250> A_IWL<17249> A_IWL<17248> A_IWL<17247> A_IWL<17246> A_IWL<17245> A_IWL<17244> A_IWL<17243> A_IWL<17242> A_IWL<17241> A_IWL<17240> A_IWL<17239> A_IWL<17238> A_IWL<17237> A_IWL<17236> A_IWL<17235> A_IWL<17234> A_IWL<17233> A_IWL<17232> A_IWL<17231> A_IWL<17230> A_IWL<17229> A_IWL<17228> A_IWL<17227> A_IWL<17226> A_IWL<17225> A_IWL<17224> A_IWL<17223> A_IWL<17222> A_IWL<17221> A_IWL<17220> A_IWL<17219> A_IWL<17218> A_IWL<17217> A_IWL<17216> A_IWL<17215> A_IWL<17214> A_IWL<17213> A_IWL<17212> A_IWL<17211> A_IWL<17210> A_IWL<17209> A_IWL<17208> A_IWL<17207> A_IWL<17206> A_IWL<17205> A_IWL<17204> A_IWL<17203> A_IWL<17202> A_IWL<17201> A_IWL<17200> A_IWL<17199> A_IWL<17198> A_IWL<17197> A_IWL<17196> A_IWL<17195> A_IWL<17194> A_IWL<17193> A_IWL<17192> A_IWL<17191> A_IWL<17190> A_IWL<17189> A_IWL<17188> A_IWL<17187> A_IWL<17186> A_IWL<17185> A_IWL<17184> A_IWL<17183> A_IWL<17182> A_IWL<17181> A_IWL<17180> A_IWL<17179> A_IWL<17178> A_IWL<17177> A_IWL<17176> A_IWL<17175> A_IWL<17174> A_IWL<17173> A_IWL<17172> A_IWL<17171> A_IWL<17170> A_IWL<17169> A_IWL<17168> A_IWL<17167> A_IWL<17166> A_IWL<17165> A_IWL<17164> A_IWL<17163> A_IWL<17162> A_IWL<17161> A_IWL<17160> A_IWL<17159> A_IWL<17158> A_IWL<17157> A_IWL<17156> A_IWL<17155> A_IWL<17154> A_IWL<17153> A_IWL<17152> A_IWL<17151> A_IWL<17150> A_IWL<17149> A_IWL<17148> A_IWL<17147> A_IWL<17146> A_IWL<17145> A_IWL<17144> A_IWL<17143> A_IWL<17142> A_IWL<17141> A_IWL<17140> A_IWL<17139> A_IWL<17138> A_IWL<17137> A_IWL<17136> A_IWL<17135> A_IWL<17134> A_IWL<17133> A_IWL<17132> A_IWL<17131> A_IWL<17130> A_IWL<17129> A_IWL<17128> A_IWL<17127> A_IWL<17126> A_IWL<17125> A_IWL<17124> A_IWL<17123> A_IWL<17122> A_IWL<17121> A_IWL<17120> A_IWL<17119> A_IWL<17118> A_IWL<17117> A_IWL<17116> A_IWL<17115> A_IWL<17114> A_IWL<17113> A_IWL<17112> A_IWL<17111> A_IWL<17110> A_IWL<17109> A_IWL<17108> A_IWL<17107> A_IWL<17106> A_IWL<17105> A_IWL<17104> A_IWL<17103> A_IWL<17102> A_IWL<17101> A_IWL<17100> A_IWL<17099> A_IWL<17098> A_IWL<17097> A_IWL<17096> A_IWL<17095> A_IWL<17094> A_IWL<17093> A_IWL<17092> A_IWL<17091> A_IWL<17090> A_IWL<17089> A_IWL<17088> A_IWL<17087> A_IWL<17086> A_IWL<17085> A_IWL<17084> A_IWL<17083> A_IWL<17082> A_IWL<17081> A_IWL<17080> A_IWL<17079> A_IWL<17078> A_IWL<17077> A_IWL<17076> A_IWL<17075> A_IWL<17074> A_IWL<17073> A_IWL<17072> A_IWL<17071> A_IWL<17070> A_IWL<17069> A_IWL<17068> A_IWL<17067> A_IWL<17066> A_IWL<17065> A_IWL<17064> A_IWL<17063> A_IWL<17062> A_IWL<17061> A_IWL<17060> A_IWL<17059> A_IWL<17058> A_IWL<17057> A_IWL<17056> A_IWL<17055> A_IWL<17054> A_IWL<17053> A_IWL<17052> A_IWL<17051> A_IWL<17050> A_IWL<17049> A_IWL<17048> A_IWL<17047> A_IWL<17046> A_IWL<17045> A_IWL<17044> A_IWL<17043> A_IWL<17042> A_IWL<17041> A_IWL<17040> A_IWL<17039> A_IWL<17038> A_IWL<17037> A_IWL<17036> A_IWL<17035> A_IWL<17034> A_IWL<17033> A_IWL<17032> A_IWL<17031> A_IWL<17030> A_IWL<17029> A_IWL<17028> A_IWL<17027> A_IWL<17026> A_IWL<17025> A_IWL<17024> A_IWL<17023> A_IWL<17022> A_IWL<17021> A_IWL<17020> A_IWL<17019> A_IWL<17018> A_IWL<17017> A_IWL<17016> A_IWL<17015> A_IWL<17014> A_IWL<17013> A_IWL<17012> A_IWL<17011> A_IWL<17010> A_IWL<17009> A_IWL<17008> A_IWL<17007> A_IWL<17006> A_IWL<17005> A_IWL<17004> A_IWL<17003> A_IWL<17002> A_IWL<17001> A_IWL<17000> A_IWL<16999> A_IWL<16998> A_IWL<16997> A_IWL<16996> A_IWL<16995> A_IWL<16994> A_IWL<16993> A_IWL<16992> A_IWL<16991> A_IWL<16990> A_IWL<16989> A_IWL<16988> A_IWL<16987> A_IWL<16986> A_IWL<16985> A_IWL<16984> A_IWL<16983> A_IWL<16982> A_IWL<16981> A_IWL<16980> A_IWL<16979> A_IWL<16978> A_IWL<16977> A_IWL<16976> A_IWL<16975> A_IWL<16974> A_IWL<16973> A_IWL<16972> A_IWL<16971> A_IWL<16970> A_IWL<16969> A_IWL<16968> A_IWL<16967> A_IWL<16966> A_IWL<16965> A_IWL<16964> A_IWL<16963> A_IWL<16962> A_IWL<16961> A_IWL<16960> A_IWL<16959> A_IWL<16958> A_IWL<16957> A_IWL<16956> A_IWL<16955> A_IWL<16954> A_IWL<16953> A_IWL<16952> A_IWL<16951> A_IWL<16950> A_IWL<16949> A_IWL<16948> A_IWL<16947> A_IWL<16946> A_IWL<16945> A_IWL<16944> A_IWL<16943> A_IWL<16942> A_IWL<16941> A_IWL<16940> A_IWL<16939> A_IWL<16938> A_IWL<16937> A_IWL<16936> A_IWL<16935> A_IWL<16934> A_IWL<16933> A_IWL<16932> A_IWL<16931> A_IWL<16930> A_IWL<16929> A_IWL<16928> A_IWL<16927> A_IWL<16926> A_IWL<16925> A_IWL<16924> A_IWL<16923> A_IWL<16922> A_IWL<16921> A_IWL<16920> A_IWL<16919> A_IWL<16918> A_IWL<16917> A_IWL<16916> A_IWL<16915> A_IWL<16914> A_IWL<16913> A_IWL<16912> A_IWL<16911> A_IWL<16910> A_IWL<16909> A_IWL<16908> A_IWL<16907> A_IWL<16906> A_IWL<16905> A_IWL<16904> A_IWL<16903> A_IWL<16902> A_IWL<16901> A_IWL<16900> A_IWL<16899> A_IWL<16898> A_IWL<16897> A_IWL<16896> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<32> A_BLC<65> A_BLC<64> A_BLC_TOP<65> A_BLC_TOP<64> A_BLT<65> A_BLT<64> A_BLT_TOP<65> A_BLT_TOP<64> A_IWL<16383> A_IWL<16382> A_IWL<16381> A_IWL<16380> A_IWL<16379> A_IWL<16378> A_IWL<16377> A_IWL<16376> A_IWL<16375> A_IWL<16374> A_IWL<16373> A_IWL<16372> A_IWL<16371> A_IWL<16370> A_IWL<16369> A_IWL<16368> A_IWL<16367> A_IWL<16366> A_IWL<16365> A_IWL<16364> A_IWL<16363> A_IWL<16362> A_IWL<16361> A_IWL<16360> A_IWL<16359> A_IWL<16358> A_IWL<16357> A_IWL<16356> A_IWL<16355> A_IWL<16354> A_IWL<16353> A_IWL<16352> A_IWL<16351> A_IWL<16350> A_IWL<16349> A_IWL<16348> A_IWL<16347> A_IWL<16346> A_IWL<16345> A_IWL<16344> A_IWL<16343> A_IWL<16342> A_IWL<16341> A_IWL<16340> A_IWL<16339> A_IWL<16338> A_IWL<16337> A_IWL<16336> A_IWL<16335> A_IWL<16334> A_IWL<16333> A_IWL<16332> A_IWL<16331> A_IWL<16330> A_IWL<16329> A_IWL<16328> A_IWL<16327> A_IWL<16326> A_IWL<16325> A_IWL<16324> A_IWL<16323> A_IWL<16322> A_IWL<16321> A_IWL<16320> A_IWL<16319> A_IWL<16318> A_IWL<16317> A_IWL<16316> A_IWL<16315> A_IWL<16314> A_IWL<16313> A_IWL<16312> A_IWL<16311> A_IWL<16310> A_IWL<16309> A_IWL<16308> A_IWL<16307> A_IWL<16306> A_IWL<16305> A_IWL<16304> A_IWL<16303> A_IWL<16302> A_IWL<16301> A_IWL<16300> A_IWL<16299> A_IWL<16298> A_IWL<16297> A_IWL<16296> A_IWL<16295> A_IWL<16294> A_IWL<16293> A_IWL<16292> A_IWL<16291> A_IWL<16290> A_IWL<16289> A_IWL<16288> A_IWL<16287> A_IWL<16286> A_IWL<16285> A_IWL<16284> A_IWL<16283> A_IWL<16282> A_IWL<16281> A_IWL<16280> A_IWL<16279> A_IWL<16278> A_IWL<16277> A_IWL<16276> A_IWL<16275> A_IWL<16274> A_IWL<16273> A_IWL<16272> A_IWL<16271> A_IWL<16270> A_IWL<16269> A_IWL<16268> A_IWL<16267> A_IWL<16266> A_IWL<16265> A_IWL<16264> A_IWL<16263> A_IWL<16262> A_IWL<16261> A_IWL<16260> A_IWL<16259> A_IWL<16258> A_IWL<16257> A_IWL<16256> A_IWL<16255> A_IWL<16254> A_IWL<16253> A_IWL<16252> A_IWL<16251> A_IWL<16250> A_IWL<16249> A_IWL<16248> A_IWL<16247> A_IWL<16246> A_IWL<16245> A_IWL<16244> A_IWL<16243> A_IWL<16242> A_IWL<16241> A_IWL<16240> A_IWL<16239> A_IWL<16238> A_IWL<16237> A_IWL<16236> A_IWL<16235> A_IWL<16234> A_IWL<16233> A_IWL<16232> A_IWL<16231> A_IWL<16230> A_IWL<16229> A_IWL<16228> A_IWL<16227> A_IWL<16226> A_IWL<16225> A_IWL<16224> A_IWL<16223> A_IWL<16222> A_IWL<16221> A_IWL<16220> A_IWL<16219> A_IWL<16218> A_IWL<16217> A_IWL<16216> A_IWL<16215> A_IWL<16214> A_IWL<16213> A_IWL<16212> A_IWL<16211> A_IWL<16210> A_IWL<16209> A_IWL<16208> A_IWL<16207> A_IWL<16206> A_IWL<16205> A_IWL<16204> A_IWL<16203> A_IWL<16202> A_IWL<16201> A_IWL<16200> A_IWL<16199> A_IWL<16198> A_IWL<16197> A_IWL<16196> A_IWL<16195> A_IWL<16194> A_IWL<16193> A_IWL<16192> A_IWL<16191> A_IWL<16190> A_IWL<16189> A_IWL<16188> A_IWL<16187> A_IWL<16186> A_IWL<16185> A_IWL<16184> A_IWL<16183> A_IWL<16182> A_IWL<16181> A_IWL<16180> A_IWL<16179> A_IWL<16178> A_IWL<16177> A_IWL<16176> A_IWL<16175> A_IWL<16174> A_IWL<16173> A_IWL<16172> A_IWL<16171> A_IWL<16170> A_IWL<16169> A_IWL<16168> A_IWL<16167> A_IWL<16166> A_IWL<16165> A_IWL<16164> A_IWL<16163> A_IWL<16162> A_IWL<16161> A_IWL<16160> A_IWL<16159> A_IWL<16158> A_IWL<16157> A_IWL<16156> A_IWL<16155> A_IWL<16154> A_IWL<16153> A_IWL<16152> A_IWL<16151> A_IWL<16150> A_IWL<16149> A_IWL<16148> A_IWL<16147> A_IWL<16146> A_IWL<16145> A_IWL<16144> A_IWL<16143> A_IWL<16142> A_IWL<16141> A_IWL<16140> A_IWL<16139> A_IWL<16138> A_IWL<16137> A_IWL<16136> A_IWL<16135> A_IWL<16134> A_IWL<16133> A_IWL<16132> A_IWL<16131> A_IWL<16130> A_IWL<16129> A_IWL<16128> A_IWL<16127> A_IWL<16126> A_IWL<16125> A_IWL<16124> A_IWL<16123> A_IWL<16122> A_IWL<16121> A_IWL<16120> A_IWL<16119> A_IWL<16118> A_IWL<16117> A_IWL<16116> A_IWL<16115> A_IWL<16114> A_IWL<16113> A_IWL<16112> A_IWL<16111> A_IWL<16110> A_IWL<16109> A_IWL<16108> A_IWL<16107> A_IWL<16106> A_IWL<16105> A_IWL<16104> A_IWL<16103> A_IWL<16102> A_IWL<16101> A_IWL<16100> A_IWL<16099> A_IWL<16098> A_IWL<16097> A_IWL<16096> A_IWL<16095> A_IWL<16094> A_IWL<16093> A_IWL<16092> A_IWL<16091> A_IWL<16090> A_IWL<16089> A_IWL<16088> A_IWL<16087> A_IWL<16086> A_IWL<16085> A_IWL<16084> A_IWL<16083> A_IWL<16082> A_IWL<16081> A_IWL<16080> A_IWL<16079> A_IWL<16078> A_IWL<16077> A_IWL<16076> A_IWL<16075> A_IWL<16074> A_IWL<16073> A_IWL<16072> A_IWL<16071> A_IWL<16070> A_IWL<16069> A_IWL<16068> A_IWL<16067> A_IWL<16066> A_IWL<16065> A_IWL<16064> A_IWL<16063> A_IWL<16062> A_IWL<16061> A_IWL<16060> A_IWL<16059> A_IWL<16058> A_IWL<16057> A_IWL<16056> A_IWL<16055> A_IWL<16054> A_IWL<16053> A_IWL<16052> A_IWL<16051> A_IWL<16050> A_IWL<16049> A_IWL<16048> A_IWL<16047> A_IWL<16046> A_IWL<16045> A_IWL<16044> A_IWL<16043> A_IWL<16042> A_IWL<16041> A_IWL<16040> A_IWL<16039> A_IWL<16038> A_IWL<16037> A_IWL<16036> A_IWL<16035> A_IWL<16034> A_IWL<16033> A_IWL<16032> A_IWL<16031> A_IWL<16030> A_IWL<16029> A_IWL<16028> A_IWL<16027> A_IWL<16026> A_IWL<16025> A_IWL<16024> A_IWL<16023> A_IWL<16022> A_IWL<16021> A_IWL<16020> A_IWL<16019> A_IWL<16018> A_IWL<16017> A_IWL<16016> A_IWL<16015> A_IWL<16014> A_IWL<16013> A_IWL<16012> A_IWL<16011> A_IWL<16010> A_IWL<16009> A_IWL<16008> A_IWL<16007> A_IWL<16006> A_IWL<16005> A_IWL<16004> A_IWL<16003> A_IWL<16002> A_IWL<16001> A_IWL<16000> A_IWL<15999> A_IWL<15998> A_IWL<15997> A_IWL<15996> A_IWL<15995> A_IWL<15994> A_IWL<15993> A_IWL<15992> A_IWL<15991> A_IWL<15990> A_IWL<15989> A_IWL<15988> A_IWL<15987> A_IWL<15986> A_IWL<15985> A_IWL<15984> A_IWL<15983> A_IWL<15982> A_IWL<15981> A_IWL<15980> A_IWL<15979> A_IWL<15978> A_IWL<15977> A_IWL<15976> A_IWL<15975> A_IWL<15974> A_IWL<15973> A_IWL<15972> A_IWL<15971> A_IWL<15970> A_IWL<15969> A_IWL<15968> A_IWL<15967> A_IWL<15966> A_IWL<15965> A_IWL<15964> A_IWL<15963> A_IWL<15962> A_IWL<15961> A_IWL<15960> A_IWL<15959> A_IWL<15958> A_IWL<15957> A_IWL<15956> A_IWL<15955> A_IWL<15954> A_IWL<15953> A_IWL<15952> A_IWL<15951> A_IWL<15950> A_IWL<15949> A_IWL<15948> A_IWL<15947> A_IWL<15946> A_IWL<15945> A_IWL<15944> A_IWL<15943> A_IWL<15942> A_IWL<15941> A_IWL<15940> A_IWL<15939> A_IWL<15938> A_IWL<15937> A_IWL<15936> A_IWL<15935> A_IWL<15934> A_IWL<15933> A_IWL<15932> A_IWL<15931> A_IWL<15930> A_IWL<15929> A_IWL<15928> A_IWL<15927> A_IWL<15926> A_IWL<15925> A_IWL<15924> A_IWL<15923> A_IWL<15922> A_IWL<15921> A_IWL<15920> A_IWL<15919> A_IWL<15918> A_IWL<15917> A_IWL<15916> A_IWL<15915> A_IWL<15914> A_IWL<15913> A_IWL<15912> A_IWL<15911> A_IWL<15910> A_IWL<15909> A_IWL<15908> A_IWL<15907> A_IWL<15906> A_IWL<15905> A_IWL<15904> A_IWL<15903> A_IWL<15902> A_IWL<15901> A_IWL<15900> A_IWL<15899> A_IWL<15898> A_IWL<15897> A_IWL<15896> A_IWL<15895> A_IWL<15894> A_IWL<15893> A_IWL<15892> A_IWL<15891> A_IWL<15890> A_IWL<15889> A_IWL<15888> A_IWL<15887> A_IWL<15886> A_IWL<15885> A_IWL<15884> A_IWL<15883> A_IWL<15882> A_IWL<15881> A_IWL<15880> A_IWL<15879> A_IWL<15878> A_IWL<15877> A_IWL<15876> A_IWL<15875> A_IWL<15874> A_IWL<15873> A_IWL<15872> A_IWL<16895> A_IWL<16894> A_IWL<16893> A_IWL<16892> A_IWL<16891> A_IWL<16890> A_IWL<16889> A_IWL<16888> A_IWL<16887> A_IWL<16886> A_IWL<16885> A_IWL<16884> A_IWL<16883> A_IWL<16882> A_IWL<16881> A_IWL<16880> A_IWL<16879> A_IWL<16878> A_IWL<16877> A_IWL<16876> A_IWL<16875> A_IWL<16874> A_IWL<16873> A_IWL<16872> A_IWL<16871> A_IWL<16870> A_IWL<16869> A_IWL<16868> A_IWL<16867> A_IWL<16866> A_IWL<16865> A_IWL<16864> A_IWL<16863> A_IWL<16862> A_IWL<16861> A_IWL<16860> A_IWL<16859> A_IWL<16858> A_IWL<16857> A_IWL<16856> A_IWL<16855> A_IWL<16854> A_IWL<16853> A_IWL<16852> A_IWL<16851> A_IWL<16850> A_IWL<16849> A_IWL<16848> A_IWL<16847> A_IWL<16846> A_IWL<16845> A_IWL<16844> A_IWL<16843> A_IWL<16842> A_IWL<16841> A_IWL<16840> A_IWL<16839> A_IWL<16838> A_IWL<16837> A_IWL<16836> A_IWL<16835> A_IWL<16834> A_IWL<16833> A_IWL<16832> A_IWL<16831> A_IWL<16830> A_IWL<16829> A_IWL<16828> A_IWL<16827> A_IWL<16826> A_IWL<16825> A_IWL<16824> A_IWL<16823> A_IWL<16822> A_IWL<16821> A_IWL<16820> A_IWL<16819> A_IWL<16818> A_IWL<16817> A_IWL<16816> A_IWL<16815> A_IWL<16814> A_IWL<16813> A_IWL<16812> A_IWL<16811> A_IWL<16810> A_IWL<16809> A_IWL<16808> A_IWL<16807> A_IWL<16806> A_IWL<16805> A_IWL<16804> A_IWL<16803> A_IWL<16802> A_IWL<16801> A_IWL<16800> A_IWL<16799> A_IWL<16798> A_IWL<16797> A_IWL<16796> A_IWL<16795> A_IWL<16794> A_IWL<16793> A_IWL<16792> A_IWL<16791> A_IWL<16790> A_IWL<16789> A_IWL<16788> A_IWL<16787> A_IWL<16786> A_IWL<16785> A_IWL<16784> A_IWL<16783> A_IWL<16782> A_IWL<16781> A_IWL<16780> A_IWL<16779> A_IWL<16778> A_IWL<16777> A_IWL<16776> A_IWL<16775> A_IWL<16774> A_IWL<16773> A_IWL<16772> A_IWL<16771> A_IWL<16770> A_IWL<16769> A_IWL<16768> A_IWL<16767> A_IWL<16766> A_IWL<16765> A_IWL<16764> A_IWL<16763> A_IWL<16762> A_IWL<16761> A_IWL<16760> A_IWL<16759> A_IWL<16758> A_IWL<16757> A_IWL<16756> A_IWL<16755> A_IWL<16754> A_IWL<16753> A_IWL<16752> A_IWL<16751> A_IWL<16750> A_IWL<16749> A_IWL<16748> A_IWL<16747> A_IWL<16746> A_IWL<16745> A_IWL<16744> A_IWL<16743> A_IWL<16742> A_IWL<16741> A_IWL<16740> A_IWL<16739> A_IWL<16738> A_IWL<16737> A_IWL<16736> A_IWL<16735> A_IWL<16734> A_IWL<16733> A_IWL<16732> A_IWL<16731> A_IWL<16730> A_IWL<16729> A_IWL<16728> A_IWL<16727> A_IWL<16726> A_IWL<16725> A_IWL<16724> A_IWL<16723> A_IWL<16722> A_IWL<16721> A_IWL<16720> A_IWL<16719> A_IWL<16718> A_IWL<16717> A_IWL<16716> A_IWL<16715> A_IWL<16714> A_IWL<16713> A_IWL<16712> A_IWL<16711> A_IWL<16710> A_IWL<16709> A_IWL<16708> A_IWL<16707> A_IWL<16706> A_IWL<16705> A_IWL<16704> A_IWL<16703> A_IWL<16702> A_IWL<16701> A_IWL<16700> A_IWL<16699> A_IWL<16698> A_IWL<16697> A_IWL<16696> A_IWL<16695> A_IWL<16694> A_IWL<16693> A_IWL<16692> A_IWL<16691> A_IWL<16690> A_IWL<16689> A_IWL<16688> A_IWL<16687> A_IWL<16686> A_IWL<16685> A_IWL<16684> A_IWL<16683> A_IWL<16682> A_IWL<16681> A_IWL<16680> A_IWL<16679> A_IWL<16678> A_IWL<16677> A_IWL<16676> A_IWL<16675> A_IWL<16674> A_IWL<16673> A_IWL<16672> A_IWL<16671> A_IWL<16670> A_IWL<16669> A_IWL<16668> A_IWL<16667> A_IWL<16666> A_IWL<16665> A_IWL<16664> A_IWL<16663> A_IWL<16662> A_IWL<16661> A_IWL<16660> A_IWL<16659> A_IWL<16658> A_IWL<16657> A_IWL<16656> A_IWL<16655> A_IWL<16654> A_IWL<16653> A_IWL<16652> A_IWL<16651> A_IWL<16650> A_IWL<16649> A_IWL<16648> A_IWL<16647> A_IWL<16646> A_IWL<16645> A_IWL<16644> A_IWL<16643> A_IWL<16642> A_IWL<16641> A_IWL<16640> A_IWL<16639> A_IWL<16638> A_IWL<16637> A_IWL<16636> A_IWL<16635> A_IWL<16634> A_IWL<16633> A_IWL<16632> A_IWL<16631> A_IWL<16630> A_IWL<16629> A_IWL<16628> A_IWL<16627> A_IWL<16626> A_IWL<16625> A_IWL<16624> A_IWL<16623> A_IWL<16622> A_IWL<16621> A_IWL<16620> A_IWL<16619> A_IWL<16618> A_IWL<16617> A_IWL<16616> A_IWL<16615> A_IWL<16614> A_IWL<16613> A_IWL<16612> A_IWL<16611> A_IWL<16610> A_IWL<16609> A_IWL<16608> A_IWL<16607> A_IWL<16606> A_IWL<16605> A_IWL<16604> A_IWL<16603> A_IWL<16602> A_IWL<16601> A_IWL<16600> A_IWL<16599> A_IWL<16598> A_IWL<16597> A_IWL<16596> A_IWL<16595> A_IWL<16594> A_IWL<16593> A_IWL<16592> A_IWL<16591> A_IWL<16590> A_IWL<16589> A_IWL<16588> A_IWL<16587> A_IWL<16586> A_IWL<16585> A_IWL<16584> A_IWL<16583> A_IWL<16582> A_IWL<16581> A_IWL<16580> A_IWL<16579> A_IWL<16578> A_IWL<16577> A_IWL<16576> A_IWL<16575> A_IWL<16574> A_IWL<16573> A_IWL<16572> A_IWL<16571> A_IWL<16570> A_IWL<16569> A_IWL<16568> A_IWL<16567> A_IWL<16566> A_IWL<16565> A_IWL<16564> A_IWL<16563> A_IWL<16562> A_IWL<16561> A_IWL<16560> A_IWL<16559> A_IWL<16558> A_IWL<16557> A_IWL<16556> A_IWL<16555> A_IWL<16554> A_IWL<16553> A_IWL<16552> A_IWL<16551> A_IWL<16550> A_IWL<16549> A_IWL<16548> A_IWL<16547> A_IWL<16546> A_IWL<16545> A_IWL<16544> A_IWL<16543> A_IWL<16542> A_IWL<16541> A_IWL<16540> A_IWL<16539> A_IWL<16538> A_IWL<16537> A_IWL<16536> A_IWL<16535> A_IWL<16534> A_IWL<16533> A_IWL<16532> A_IWL<16531> A_IWL<16530> A_IWL<16529> A_IWL<16528> A_IWL<16527> A_IWL<16526> A_IWL<16525> A_IWL<16524> A_IWL<16523> A_IWL<16522> A_IWL<16521> A_IWL<16520> A_IWL<16519> A_IWL<16518> A_IWL<16517> A_IWL<16516> A_IWL<16515> A_IWL<16514> A_IWL<16513> A_IWL<16512> A_IWL<16511> A_IWL<16510> A_IWL<16509> A_IWL<16508> A_IWL<16507> A_IWL<16506> A_IWL<16505> A_IWL<16504> A_IWL<16503> A_IWL<16502> A_IWL<16501> A_IWL<16500> A_IWL<16499> A_IWL<16498> A_IWL<16497> A_IWL<16496> A_IWL<16495> A_IWL<16494> A_IWL<16493> A_IWL<16492> A_IWL<16491> A_IWL<16490> A_IWL<16489> A_IWL<16488> A_IWL<16487> A_IWL<16486> A_IWL<16485> A_IWL<16484> A_IWL<16483> A_IWL<16482> A_IWL<16481> A_IWL<16480> A_IWL<16479> A_IWL<16478> A_IWL<16477> A_IWL<16476> A_IWL<16475> A_IWL<16474> A_IWL<16473> A_IWL<16472> A_IWL<16471> A_IWL<16470> A_IWL<16469> A_IWL<16468> A_IWL<16467> A_IWL<16466> A_IWL<16465> A_IWL<16464> A_IWL<16463> A_IWL<16462> A_IWL<16461> A_IWL<16460> A_IWL<16459> A_IWL<16458> A_IWL<16457> A_IWL<16456> A_IWL<16455> A_IWL<16454> A_IWL<16453> A_IWL<16452> A_IWL<16451> A_IWL<16450> A_IWL<16449> A_IWL<16448> A_IWL<16447> A_IWL<16446> A_IWL<16445> A_IWL<16444> A_IWL<16443> A_IWL<16442> A_IWL<16441> A_IWL<16440> A_IWL<16439> A_IWL<16438> A_IWL<16437> A_IWL<16436> A_IWL<16435> A_IWL<16434> A_IWL<16433> A_IWL<16432> A_IWL<16431> A_IWL<16430> A_IWL<16429> A_IWL<16428> A_IWL<16427> A_IWL<16426> A_IWL<16425> A_IWL<16424> A_IWL<16423> A_IWL<16422> A_IWL<16421> A_IWL<16420> A_IWL<16419> A_IWL<16418> A_IWL<16417> A_IWL<16416> A_IWL<16415> A_IWL<16414> A_IWL<16413> A_IWL<16412> A_IWL<16411> A_IWL<16410> A_IWL<16409> A_IWL<16408> A_IWL<16407> A_IWL<16406> A_IWL<16405> A_IWL<16404> A_IWL<16403> A_IWL<16402> A_IWL<16401> A_IWL<16400> A_IWL<16399> A_IWL<16398> A_IWL<16397> A_IWL<16396> A_IWL<16395> A_IWL<16394> A_IWL<16393> A_IWL<16392> A_IWL<16391> A_IWL<16390> A_IWL<16389> A_IWL<16388> A_IWL<16387> A_IWL<16386> A_IWL<16385> A_IWL<16384> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<31> A_BLC<63> A_BLC<62> A_BLC_TOP<63> A_BLC_TOP<62> A_BLT<63> A_BLT<62> A_BLT_TOP<63> A_BLT_TOP<62> A_IWL<15871> A_IWL<15870> A_IWL<15869> A_IWL<15868> A_IWL<15867> A_IWL<15866> A_IWL<15865> A_IWL<15864> A_IWL<15863> A_IWL<15862> A_IWL<15861> A_IWL<15860> A_IWL<15859> A_IWL<15858> A_IWL<15857> A_IWL<15856> A_IWL<15855> A_IWL<15854> A_IWL<15853> A_IWL<15852> A_IWL<15851> A_IWL<15850> A_IWL<15849> A_IWL<15848> A_IWL<15847> A_IWL<15846> A_IWL<15845> A_IWL<15844> A_IWL<15843> A_IWL<15842> A_IWL<15841> A_IWL<15840> A_IWL<15839> A_IWL<15838> A_IWL<15837> A_IWL<15836> A_IWL<15835> A_IWL<15834> A_IWL<15833> A_IWL<15832> A_IWL<15831> A_IWL<15830> A_IWL<15829> A_IWL<15828> A_IWL<15827> A_IWL<15826> A_IWL<15825> A_IWL<15824> A_IWL<15823> A_IWL<15822> A_IWL<15821> A_IWL<15820> A_IWL<15819> A_IWL<15818> A_IWL<15817> A_IWL<15816> A_IWL<15815> A_IWL<15814> A_IWL<15813> A_IWL<15812> A_IWL<15811> A_IWL<15810> A_IWL<15809> A_IWL<15808> A_IWL<15807> A_IWL<15806> A_IWL<15805> A_IWL<15804> A_IWL<15803> A_IWL<15802> A_IWL<15801> A_IWL<15800> A_IWL<15799> A_IWL<15798> A_IWL<15797> A_IWL<15796> A_IWL<15795> A_IWL<15794> A_IWL<15793> A_IWL<15792> A_IWL<15791> A_IWL<15790> A_IWL<15789> A_IWL<15788> A_IWL<15787> A_IWL<15786> A_IWL<15785> A_IWL<15784> A_IWL<15783> A_IWL<15782> A_IWL<15781> A_IWL<15780> A_IWL<15779> A_IWL<15778> A_IWL<15777> A_IWL<15776> A_IWL<15775> A_IWL<15774> A_IWL<15773> A_IWL<15772> A_IWL<15771> A_IWL<15770> A_IWL<15769> A_IWL<15768> A_IWL<15767> A_IWL<15766> A_IWL<15765> A_IWL<15764> A_IWL<15763> A_IWL<15762> A_IWL<15761> A_IWL<15760> A_IWL<15759> A_IWL<15758> A_IWL<15757> A_IWL<15756> A_IWL<15755> A_IWL<15754> A_IWL<15753> A_IWL<15752> A_IWL<15751> A_IWL<15750> A_IWL<15749> A_IWL<15748> A_IWL<15747> A_IWL<15746> A_IWL<15745> A_IWL<15744> A_IWL<15743> A_IWL<15742> A_IWL<15741> A_IWL<15740> A_IWL<15739> A_IWL<15738> A_IWL<15737> A_IWL<15736> A_IWL<15735> A_IWL<15734> A_IWL<15733> A_IWL<15732> A_IWL<15731> A_IWL<15730> A_IWL<15729> A_IWL<15728> A_IWL<15727> A_IWL<15726> A_IWL<15725> A_IWL<15724> A_IWL<15723> A_IWL<15722> A_IWL<15721> A_IWL<15720> A_IWL<15719> A_IWL<15718> A_IWL<15717> A_IWL<15716> A_IWL<15715> A_IWL<15714> A_IWL<15713> A_IWL<15712> A_IWL<15711> A_IWL<15710> A_IWL<15709> A_IWL<15708> A_IWL<15707> A_IWL<15706> A_IWL<15705> A_IWL<15704> A_IWL<15703> A_IWL<15702> A_IWL<15701> A_IWL<15700> A_IWL<15699> A_IWL<15698> A_IWL<15697> A_IWL<15696> A_IWL<15695> A_IWL<15694> A_IWL<15693> A_IWL<15692> A_IWL<15691> A_IWL<15690> A_IWL<15689> A_IWL<15688> A_IWL<15687> A_IWL<15686> A_IWL<15685> A_IWL<15684> A_IWL<15683> A_IWL<15682> A_IWL<15681> A_IWL<15680> A_IWL<15679> A_IWL<15678> A_IWL<15677> A_IWL<15676> A_IWL<15675> A_IWL<15674> A_IWL<15673> A_IWL<15672> A_IWL<15671> A_IWL<15670> A_IWL<15669> A_IWL<15668> A_IWL<15667> A_IWL<15666> A_IWL<15665> A_IWL<15664> A_IWL<15663> A_IWL<15662> A_IWL<15661> A_IWL<15660> A_IWL<15659> A_IWL<15658> A_IWL<15657> A_IWL<15656> A_IWL<15655> A_IWL<15654> A_IWL<15653> A_IWL<15652> A_IWL<15651> A_IWL<15650> A_IWL<15649> A_IWL<15648> A_IWL<15647> A_IWL<15646> A_IWL<15645> A_IWL<15644> A_IWL<15643> A_IWL<15642> A_IWL<15641> A_IWL<15640> A_IWL<15639> A_IWL<15638> A_IWL<15637> A_IWL<15636> A_IWL<15635> A_IWL<15634> A_IWL<15633> A_IWL<15632> A_IWL<15631> A_IWL<15630> A_IWL<15629> A_IWL<15628> A_IWL<15627> A_IWL<15626> A_IWL<15625> A_IWL<15624> A_IWL<15623> A_IWL<15622> A_IWL<15621> A_IWL<15620> A_IWL<15619> A_IWL<15618> A_IWL<15617> A_IWL<15616> A_IWL<15615> A_IWL<15614> A_IWL<15613> A_IWL<15612> A_IWL<15611> A_IWL<15610> A_IWL<15609> A_IWL<15608> A_IWL<15607> A_IWL<15606> A_IWL<15605> A_IWL<15604> A_IWL<15603> A_IWL<15602> A_IWL<15601> A_IWL<15600> A_IWL<15599> A_IWL<15598> A_IWL<15597> A_IWL<15596> A_IWL<15595> A_IWL<15594> A_IWL<15593> A_IWL<15592> A_IWL<15591> A_IWL<15590> A_IWL<15589> A_IWL<15588> A_IWL<15587> A_IWL<15586> A_IWL<15585> A_IWL<15584> A_IWL<15583> A_IWL<15582> A_IWL<15581> A_IWL<15580> A_IWL<15579> A_IWL<15578> A_IWL<15577> A_IWL<15576> A_IWL<15575> A_IWL<15574> A_IWL<15573> A_IWL<15572> A_IWL<15571> A_IWL<15570> A_IWL<15569> A_IWL<15568> A_IWL<15567> A_IWL<15566> A_IWL<15565> A_IWL<15564> A_IWL<15563> A_IWL<15562> A_IWL<15561> A_IWL<15560> A_IWL<15559> A_IWL<15558> A_IWL<15557> A_IWL<15556> A_IWL<15555> A_IWL<15554> A_IWL<15553> A_IWL<15552> A_IWL<15551> A_IWL<15550> A_IWL<15549> A_IWL<15548> A_IWL<15547> A_IWL<15546> A_IWL<15545> A_IWL<15544> A_IWL<15543> A_IWL<15542> A_IWL<15541> A_IWL<15540> A_IWL<15539> A_IWL<15538> A_IWL<15537> A_IWL<15536> A_IWL<15535> A_IWL<15534> A_IWL<15533> A_IWL<15532> A_IWL<15531> A_IWL<15530> A_IWL<15529> A_IWL<15528> A_IWL<15527> A_IWL<15526> A_IWL<15525> A_IWL<15524> A_IWL<15523> A_IWL<15522> A_IWL<15521> A_IWL<15520> A_IWL<15519> A_IWL<15518> A_IWL<15517> A_IWL<15516> A_IWL<15515> A_IWL<15514> A_IWL<15513> A_IWL<15512> A_IWL<15511> A_IWL<15510> A_IWL<15509> A_IWL<15508> A_IWL<15507> A_IWL<15506> A_IWL<15505> A_IWL<15504> A_IWL<15503> A_IWL<15502> A_IWL<15501> A_IWL<15500> A_IWL<15499> A_IWL<15498> A_IWL<15497> A_IWL<15496> A_IWL<15495> A_IWL<15494> A_IWL<15493> A_IWL<15492> A_IWL<15491> A_IWL<15490> A_IWL<15489> A_IWL<15488> A_IWL<15487> A_IWL<15486> A_IWL<15485> A_IWL<15484> A_IWL<15483> A_IWL<15482> A_IWL<15481> A_IWL<15480> A_IWL<15479> A_IWL<15478> A_IWL<15477> A_IWL<15476> A_IWL<15475> A_IWL<15474> A_IWL<15473> A_IWL<15472> A_IWL<15471> A_IWL<15470> A_IWL<15469> A_IWL<15468> A_IWL<15467> A_IWL<15466> A_IWL<15465> A_IWL<15464> A_IWL<15463> A_IWL<15462> A_IWL<15461> A_IWL<15460> A_IWL<15459> A_IWL<15458> A_IWL<15457> A_IWL<15456> A_IWL<15455> A_IWL<15454> A_IWL<15453> A_IWL<15452> A_IWL<15451> A_IWL<15450> A_IWL<15449> A_IWL<15448> A_IWL<15447> A_IWL<15446> A_IWL<15445> A_IWL<15444> A_IWL<15443> A_IWL<15442> A_IWL<15441> A_IWL<15440> A_IWL<15439> A_IWL<15438> A_IWL<15437> A_IWL<15436> A_IWL<15435> A_IWL<15434> A_IWL<15433> A_IWL<15432> A_IWL<15431> A_IWL<15430> A_IWL<15429> A_IWL<15428> A_IWL<15427> A_IWL<15426> A_IWL<15425> A_IWL<15424> A_IWL<15423> A_IWL<15422> A_IWL<15421> A_IWL<15420> A_IWL<15419> A_IWL<15418> A_IWL<15417> A_IWL<15416> A_IWL<15415> A_IWL<15414> A_IWL<15413> A_IWL<15412> A_IWL<15411> A_IWL<15410> A_IWL<15409> A_IWL<15408> A_IWL<15407> A_IWL<15406> A_IWL<15405> A_IWL<15404> A_IWL<15403> A_IWL<15402> A_IWL<15401> A_IWL<15400> A_IWL<15399> A_IWL<15398> A_IWL<15397> A_IWL<15396> A_IWL<15395> A_IWL<15394> A_IWL<15393> A_IWL<15392> A_IWL<15391> A_IWL<15390> A_IWL<15389> A_IWL<15388> A_IWL<15387> A_IWL<15386> A_IWL<15385> A_IWL<15384> A_IWL<15383> A_IWL<15382> A_IWL<15381> A_IWL<15380> A_IWL<15379> A_IWL<15378> A_IWL<15377> A_IWL<15376> A_IWL<15375> A_IWL<15374> A_IWL<15373> A_IWL<15372> A_IWL<15371> A_IWL<15370> A_IWL<15369> A_IWL<15368> A_IWL<15367> A_IWL<15366> A_IWL<15365> A_IWL<15364> A_IWL<15363> A_IWL<15362> A_IWL<15361> A_IWL<15360> A_IWL<16383> A_IWL<16382> A_IWL<16381> A_IWL<16380> A_IWL<16379> A_IWL<16378> A_IWL<16377> A_IWL<16376> A_IWL<16375> A_IWL<16374> A_IWL<16373> A_IWL<16372> A_IWL<16371> A_IWL<16370> A_IWL<16369> A_IWL<16368> A_IWL<16367> A_IWL<16366> A_IWL<16365> A_IWL<16364> A_IWL<16363> A_IWL<16362> A_IWL<16361> A_IWL<16360> A_IWL<16359> A_IWL<16358> A_IWL<16357> A_IWL<16356> A_IWL<16355> A_IWL<16354> A_IWL<16353> A_IWL<16352> A_IWL<16351> A_IWL<16350> A_IWL<16349> A_IWL<16348> A_IWL<16347> A_IWL<16346> A_IWL<16345> A_IWL<16344> A_IWL<16343> A_IWL<16342> A_IWL<16341> A_IWL<16340> A_IWL<16339> A_IWL<16338> A_IWL<16337> A_IWL<16336> A_IWL<16335> A_IWL<16334> A_IWL<16333> A_IWL<16332> A_IWL<16331> A_IWL<16330> A_IWL<16329> A_IWL<16328> A_IWL<16327> A_IWL<16326> A_IWL<16325> A_IWL<16324> A_IWL<16323> A_IWL<16322> A_IWL<16321> A_IWL<16320> A_IWL<16319> A_IWL<16318> A_IWL<16317> A_IWL<16316> A_IWL<16315> A_IWL<16314> A_IWL<16313> A_IWL<16312> A_IWL<16311> A_IWL<16310> A_IWL<16309> A_IWL<16308> A_IWL<16307> A_IWL<16306> A_IWL<16305> A_IWL<16304> A_IWL<16303> A_IWL<16302> A_IWL<16301> A_IWL<16300> A_IWL<16299> A_IWL<16298> A_IWL<16297> A_IWL<16296> A_IWL<16295> A_IWL<16294> A_IWL<16293> A_IWL<16292> A_IWL<16291> A_IWL<16290> A_IWL<16289> A_IWL<16288> A_IWL<16287> A_IWL<16286> A_IWL<16285> A_IWL<16284> A_IWL<16283> A_IWL<16282> A_IWL<16281> A_IWL<16280> A_IWL<16279> A_IWL<16278> A_IWL<16277> A_IWL<16276> A_IWL<16275> A_IWL<16274> A_IWL<16273> A_IWL<16272> A_IWL<16271> A_IWL<16270> A_IWL<16269> A_IWL<16268> A_IWL<16267> A_IWL<16266> A_IWL<16265> A_IWL<16264> A_IWL<16263> A_IWL<16262> A_IWL<16261> A_IWL<16260> A_IWL<16259> A_IWL<16258> A_IWL<16257> A_IWL<16256> A_IWL<16255> A_IWL<16254> A_IWL<16253> A_IWL<16252> A_IWL<16251> A_IWL<16250> A_IWL<16249> A_IWL<16248> A_IWL<16247> A_IWL<16246> A_IWL<16245> A_IWL<16244> A_IWL<16243> A_IWL<16242> A_IWL<16241> A_IWL<16240> A_IWL<16239> A_IWL<16238> A_IWL<16237> A_IWL<16236> A_IWL<16235> A_IWL<16234> A_IWL<16233> A_IWL<16232> A_IWL<16231> A_IWL<16230> A_IWL<16229> A_IWL<16228> A_IWL<16227> A_IWL<16226> A_IWL<16225> A_IWL<16224> A_IWL<16223> A_IWL<16222> A_IWL<16221> A_IWL<16220> A_IWL<16219> A_IWL<16218> A_IWL<16217> A_IWL<16216> A_IWL<16215> A_IWL<16214> A_IWL<16213> A_IWL<16212> A_IWL<16211> A_IWL<16210> A_IWL<16209> A_IWL<16208> A_IWL<16207> A_IWL<16206> A_IWL<16205> A_IWL<16204> A_IWL<16203> A_IWL<16202> A_IWL<16201> A_IWL<16200> A_IWL<16199> A_IWL<16198> A_IWL<16197> A_IWL<16196> A_IWL<16195> A_IWL<16194> A_IWL<16193> A_IWL<16192> A_IWL<16191> A_IWL<16190> A_IWL<16189> A_IWL<16188> A_IWL<16187> A_IWL<16186> A_IWL<16185> A_IWL<16184> A_IWL<16183> A_IWL<16182> A_IWL<16181> A_IWL<16180> A_IWL<16179> A_IWL<16178> A_IWL<16177> A_IWL<16176> A_IWL<16175> A_IWL<16174> A_IWL<16173> A_IWL<16172> A_IWL<16171> A_IWL<16170> A_IWL<16169> A_IWL<16168> A_IWL<16167> A_IWL<16166> A_IWL<16165> A_IWL<16164> A_IWL<16163> A_IWL<16162> A_IWL<16161> A_IWL<16160> A_IWL<16159> A_IWL<16158> A_IWL<16157> A_IWL<16156> A_IWL<16155> A_IWL<16154> A_IWL<16153> A_IWL<16152> A_IWL<16151> A_IWL<16150> A_IWL<16149> A_IWL<16148> A_IWL<16147> A_IWL<16146> A_IWL<16145> A_IWL<16144> A_IWL<16143> A_IWL<16142> A_IWL<16141> A_IWL<16140> A_IWL<16139> A_IWL<16138> A_IWL<16137> A_IWL<16136> A_IWL<16135> A_IWL<16134> A_IWL<16133> A_IWL<16132> A_IWL<16131> A_IWL<16130> A_IWL<16129> A_IWL<16128> A_IWL<16127> A_IWL<16126> A_IWL<16125> A_IWL<16124> A_IWL<16123> A_IWL<16122> A_IWL<16121> A_IWL<16120> A_IWL<16119> A_IWL<16118> A_IWL<16117> A_IWL<16116> A_IWL<16115> A_IWL<16114> A_IWL<16113> A_IWL<16112> A_IWL<16111> A_IWL<16110> A_IWL<16109> A_IWL<16108> A_IWL<16107> A_IWL<16106> A_IWL<16105> A_IWL<16104> A_IWL<16103> A_IWL<16102> A_IWL<16101> A_IWL<16100> A_IWL<16099> A_IWL<16098> A_IWL<16097> A_IWL<16096> A_IWL<16095> A_IWL<16094> A_IWL<16093> A_IWL<16092> A_IWL<16091> A_IWL<16090> A_IWL<16089> A_IWL<16088> A_IWL<16087> A_IWL<16086> A_IWL<16085> A_IWL<16084> A_IWL<16083> A_IWL<16082> A_IWL<16081> A_IWL<16080> A_IWL<16079> A_IWL<16078> A_IWL<16077> A_IWL<16076> A_IWL<16075> A_IWL<16074> A_IWL<16073> A_IWL<16072> A_IWL<16071> A_IWL<16070> A_IWL<16069> A_IWL<16068> A_IWL<16067> A_IWL<16066> A_IWL<16065> A_IWL<16064> A_IWL<16063> A_IWL<16062> A_IWL<16061> A_IWL<16060> A_IWL<16059> A_IWL<16058> A_IWL<16057> A_IWL<16056> A_IWL<16055> A_IWL<16054> A_IWL<16053> A_IWL<16052> A_IWL<16051> A_IWL<16050> A_IWL<16049> A_IWL<16048> A_IWL<16047> A_IWL<16046> A_IWL<16045> A_IWL<16044> A_IWL<16043> A_IWL<16042> A_IWL<16041> A_IWL<16040> A_IWL<16039> A_IWL<16038> A_IWL<16037> A_IWL<16036> A_IWL<16035> A_IWL<16034> A_IWL<16033> A_IWL<16032> A_IWL<16031> A_IWL<16030> A_IWL<16029> A_IWL<16028> A_IWL<16027> A_IWL<16026> A_IWL<16025> A_IWL<16024> A_IWL<16023> A_IWL<16022> A_IWL<16021> A_IWL<16020> A_IWL<16019> A_IWL<16018> A_IWL<16017> A_IWL<16016> A_IWL<16015> A_IWL<16014> A_IWL<16013> A_IWL<16012> A_IWL<16011> A_IWL<16010> A_IWL<16009> A_IWL<16008> A_IWL<16007> A_IWL<16006> A_IWL<16005> A_IWL<16004> A_IWL<16003> A_IWL<16002> A_IWL<16001> A_IWL<16000> A_IWL<15999> A_IWL<15998> A_IWL<15997> A_IWL<15996> A_IWL<15995> A_IWL<15994> A_IWL<15993> A_IWL<15992> A_IWL<15991> A_IWL<15990> A_IWL<15989> A_IWL<15988> A_IWL<15987> A_IWL<15986> A_IWL<15985> A_IWL<15984> A_IWL<15983> A_IWL<15982> A_IWL<15981> A_IWL<15980> A_IWL<15979> A_IWL<15978> A_IWL<15977> A_IWL<15976> A_IWL<15975> A_IWL<15974> A_IWL<15973> A_IWL<15972> A_IWL<15971> A_IWL<15970> A_IWL<15969> A_IWL<15968> A_IWL<15967> A_IWL<15966> A_IWL<15965> A_IWL<15964> A_IWL<15963> A_IWL<15962> A_IWL<15961> A_IWL<15960> A_IWL<15959> A_IWL<15958> A_IWL<15957> A_IWL<15956> A_IWL<15955> A_IWL<15954> A_IWL<15953> A_IWL<15952> A_IWL<15951> A_IWL<15950> A_IWL<15949> A_IWL<15948> A_IWL<15947> A_IWL<15946> A_IWL<15945> A_IWL<15944> A_IWL<15943> A_IWL<15942> A_IWL<15941> A_IWL<15940> A_IWL<15939> A_IWL<15938> A_IWL<15937> A_IWL<15936> A_IWL<15935> A_IWL<15934> A_IWL<15933> A_IWL<15932> A_IWL<15931> A_IWL<15930> A_IWL<15929> A_IWL<15928> A_IWL<15927> A_IWL<15926> A_IWL<15925> A_IWL<15924> A_IWL<15923> A_IWL<15922> A_IWL<15921> A_IWL<15920> A_IWL<15919> A_IWL<15918> A_IWL<15917> A_IWL<15916> A_IWL<15915> A_IWL<15914> A_IWL<15913> A_IWL<15912> A_IWL<15911> A_IWL<15910> A_IWL<15909> A_IWL<15908> A_IWL<15907> A_IWL<15906> A_IWL<15905> A_IWL<15904> A_IWL<15903> A_IWL<15902> A_IWL<15901> A_IWL<15900> A_IWL<15899> A_IWL<15898> A_IWL<15897> A_IWL<15896> A_IWL<15895> A_IWL<15894> A_IWL<15893> A_IWL<15892> A_IWL<15891> A_IWL<15890> A_IWL<15889> A_IWL<15888> A_IWL<15887> A_IWL<15886> A_IWL<15885> A_IWL<15884> A_IWL<15883> A_IWL<15882> A_IWL<15881> A_IWL<15880> A_IWL<15879> A_IWL<15878> A_IWL<15877> A_IWL<15876> A_IWL<15875> A_IWL<15874> A_IWL<15873> A_IWL<15872> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<30> A_BLC<61> A_BLC<60> A_BLC_TOP<61> A_BLC_TOP<60> A_BLT<61> A_BLT<60> A_BLT_TOP<61> A_BLT_TOP<60> A_IWL<15359> A_IWL<15358> A_IWL<15357> A_IWL<15356> A_IWL<15355> A_IWL<15354> A_IWL<15353> A_IWL<15352> A_IWL<15351> A_IWL<15350> A_IWL<15349> A_IWL<15348> A_IWL<15347> A_IWL<15346> A_IWL<15345> A_IWL<15344> A_IWL<15343> A_IWL<15342> A_IWL<15341> A_IWL<15340> A_IWL<15339> A_IWL<15338> A_IWL<15337> A_IWL<15336> A_IWL<15335> A_IWL<15334> A_IWL<15333> A_IWL<15332> A_IWL<15331> A_IWL<15330> A_IWL<15329> A_IWL<15328> A_IWL<15327> A_IWL<15326> A_IWL<15325> A_IWL<15324> A_IWL<15323> A_IWL<15322> A_IWL<15321> A_IWL<15320> A_IWL<15319> A_IWL<15318> A_IWL<15317> A_IWL<15316> A_IWL<15315> A_IWL<15314> A_IWL<15313> A_IWL<15312> A_IWL<15311> A_IWL<15310> A_IWL<15309> A_IWL<15308> A_IWL<15307> A_IWL<15306> A_IWL<15305> A_IWL<15304> A_IWL<15303> A_IWL<15302> A_IWL<15301> A_IWL<15300> A_IWL<15299> A_IWL<15298> A_IWL<15297> A_IWL<15296> A_IWL<15295> A_IWL<15294> A_IWL<15293> A_IWL<15292> A_IWL<15291> A_IWL<15290> A_IWL<15289> A_IWL<15288> A_IWL<15287> A_IWL<15286> A_IWL<15285> A_IWL<15284> A_IWL<15283> A_IWL<15282> A_IWL<15281> A_IWL<15280> A_IWL<15279> A_IWL<15278> A_IWL<15277> A_IWL<15276> A_IWL<15275> A_IWL<15274> A_IWL<15273> A_IWL<15272> A_IWL<15271> A_IWL<15270> A_IWL<15269> A_IWL<15268> A_IWL<15267> A_IWL<15266> A_IWL<15265> A_IWL<15264> A_IWL<15263> A_IWL<15262> A_IWL<15261> A_IWL<15260> A_IWL<15259> A_IWL<15258> A_IWL<15257> A_IWL<15256> A_IWL<15255> A_IWL<15254> A_IWL<15253> A_IWL<15252> A_IWL<15251> A_IWL<15250> A_IWL<15249> A_IWL<15248> A_IWL<15247> A_IWL<15246> A_IWL<15245> A_IWL<15244> A_IWL<15243> A_IWL<15242> A_IWL<15241> A_IWL<15240> A_IWL<15239> A_IWL<15238> A_IWL<15237> A_IWL<15236> A_IWL<15235> A_IWL<15234> A_IWL<15233> A_IWL<15232> A_IWL<15231> A_IWL<15230> A_IWL<15229> A_IWL<15228> A_IWL<15227> A_IWL<15226> A_IWL<15225> A_IWL<15224> A_IWL<15223> A_IWL<15222> A_IWL<15221> A_IWL<15220> A_IWL<15219> A_IWL<15218> A_IWL<15217> A_IWL<15216> A_IWL<15215> A_IWL<15214> A_IWL<15213> A_IWL<15212> A_IWL<15211> A_IWL<15210> A_IWL<15209> A_IWL<15208> A_IWL<15207> A_IWL<15206> A_IWL<15205> A_IWL<15204> A_IWL<15203> A_IWL<15202> A_IWL<15201> A_IWL<15200> A_IWL<15199> A_IWL<15198> A_IWL<15197> A_IWL<15196> A_IWL<15195> A_IWL<15194> A_IWL<15193> A_IWL<15192> A_IWL<15191> A_IWL<15190> A_IWL<15189> A_IWL<15188> A_IWL<15187> A_IWL<15186> A_IWL<15185> A_IWL<15184> A_IWL<15183> A_IWL<15182> A_IWL<15181> A_IWL<15180> A_IWL<15179> A_IWL<15178> A_IWL<15177> A_IWL<15176> A_IWL<15175> A_IWL<15174> A_IWL<15173> A_IWL<15172> A_IWL<15171> A_IWL<15170> A_IWL<15169> A_IWL<15168> A_IWL<15167> A_IWL<15166> A_IWL<15165> A_IWL<15164> A_IWL<15163> A_IWL<15162> A_IWL<15161> A_IWL<15160> A_IWL<15159> A_IWL<15158> A_IWL<15157> A_IWL<15156> A_IWL<15155> A_IWL<15154> A_IWL<15153> A_IWL<15152> A_IWL<15151> A_IWL<15150> A_IWL<15149> A_IWL<15148> A_IWL<15147> A_IWL<15146> A_IWL<15145> A_IWL<15144> A_IWL<15143> A_IWL<15142> A_IWL<15141> A_IWL<15140> A_IWL<15139> A_IWL<15138> A_IWL<15137> A_IWL<15136> A_IWL<15135> A_IWL<15134> A_IWL<15133> A_IWL<15132> A_IWL<15131> A_IWL<15130> A_IWL<15129> A_IWL<15128> A_IWL<15127> A_IWL<15126> A_IWL<15125> A_IWL<15124> A_IWL<15123> A_IWL<15122> A_IWL<15121> A_IWL<15120> A_IWL<15119> A_IWL<15118> A_IWL<15117> A_IWL<15116> A_IWL<15115> A_IWL<15114> A_IWL<15113> A_IWL<15112> A_IWL<15111> A_IWL<15110> A_IWL<15109> A_IWL<15108> A_IWL<15107> A_IWL<15106> A_IWL<15105> A_IWL<15104> A_IWL<15103> A_IWL<15102> A_IWL<15101> A_IWL<15100> A_IWL<15099> A_IWL<15098> A_IWL<15097> A_IWL<15096> A_IWL<15095> A_IWL<15094> A_IWL<15093> A_IWL<15092> A_IWL<15091> A_IWL<15090> A_IWL<15089> A_IWL<15088> A_IWL<15087> A_IWL<15086> A_IWL<15085> A_IWL<15084> A_IWL<15083> A_IWL<15082> A_IWL<15081> A_IWL<15080> A_IWL<15079> A_IWL<15078> A_IWL<15077> A_IWL<15076> A_IWL<15075> A_IWL<15074> A_IWL<15073> A_IWL<15072> A_IWL<15071> A_IWL<15070> A_IWL<15069> A_IWL<15068> A_IWL<15067> A_IWL<15066> A_IWL<15065> A_IWL<15064> A_IWL<15063> A_IWL<15062> A_IWL<15061> A_IWL<15060> A_IWL<15059> A_IWL<15058> A_IWL<15057> A_IWL<15056> A_IWL<15055> A_IWL<15054> A_IWL<15053> A_IWL<15052> A_IWL<15051> A_IWL<15050> A_IWL<15049> A_IWL<15048> A_IWL<15047> A_IWL<15046> A_IWL<15045> A_IWL<15044> A_IWL<15043> A_IWL<15042> A_IWL<15041> A_IWL<15040> A_IWL<15039> A_IWL<15038> A_IWL<15037> A_IWL<15036> A_IWL<15035> A_IWL<15034> A_IWL<15033> A_IWL<15032> A_IWL<15031> A_IWL<15030> A_IWL<15029> A_IWL<15028> A_IWL<15027> A_IWL<15026> A_IWL<15025> A_IWL<15024> A_IWL<15023> A_IWL<15022> A_IWL<15021> A_IWL<15020> A_IWL<15019> A_IWL<15018> A_IWL<15017> A_IWL<15016> A_IWL<15015> A_IWL<15014> A_IWL<15013> A_IWL<15012> A_IWL<15011> A_IWL<15010> A_IWL<15009> A_IWL<15008> A_IWL<15007> A_IWL<15006> A_IWL<15005> A_IWL<15004> A_IWL<15003> A_IWL<15002> A_IWL<15001> A_IWL<15000> A_IWL<14999> A_IWL<14998> A_IWL<14997> A_IWL<14996> A_IWL<14995> A_IWL<14994> A_IWL<14993> A_IWL<14992> A_IWL<14991> A_IWL<14990> A_IWL<14989> A_IWL<14988> A_IWL<14987> A_IWL<14986> A_IWL<14985> A_IWL<14984> A_IWL<14983> A_IWL<14982> A_IWL<14981> A_IWL<14980> A_IWL<14979> A_IWL<14978> A_IWL<14977> A_IWL<14976> A_IWL<14975> A_IWL<14974> A_IWL<14973> A_IWL<14972> A_IWL<14971> A_IWL<14970> A_IWL<14969> A_IWL<14968> A_IWL<14967> A_IWL<14966> A_IWL<14965> A_IWL<14964> A_IWL<14963> A_IWL<14962> A_IWL<14961> A_IWL<14960> A_IWL<14959> A_IWL<14958> A_IWL<14957> A_IWL<14956> A_IWL<14955> A_IWL<14954> A_IWL<14953> A_IWL<14952> A_IWL<14951> A_IWL<14950> A_IWL<14949> A_IWL<14948> A_IWL<14947> A_IWL<14946> A_IWL<14945> A_IWL<14944> A_IWL<14943> A_IWL<14942> A_IWL<14941> A_IWL<14940> A_IWL<14939> A_IWL<14938> A_IWL<14937> A_IWL<14936> A_IWL<14935> A_IWL<14934> A_IWL<14933> A_IWL<14932> A_IWL<14931> A_IWL<14930> A_IWL<14929> A_IWL<14928> A_IWL<14927> A_IWL<14926> A_IWL<14925> A_IWL<14924> A_IWL<14923> A_IWL<14922> A_IWL<14921> A_IWL<14920> A_IWL<14919> A_IWL<14918> A_IWL<14917> A_IWL<14916> A_IWL<14915> A_IWL<14914> A_IWL<14913> A_IWL<14912> A_IWL<14911> A_IWL<14910> A_IWL<14909> A_IWL<14908> A_IWL<14907> A_IWL<14906> A_IWL<14905> A_IWL<14904> A_IWL<14903> A_IWL<14902> A_IWL<14901> A_IWL<14900> A_IWL<14899> A_IWL<14898> A_IWL<14897> A_IWL<14896> A_IWL<14895> A_IWL<14894> A_IWL<14893> A_IWL<14892> A_IWL<14891> A_IWL<14890> A_IWL<14889> A_IWL<14888> A_IWL<14887> A_IWL<14886> A_IWL<14885> A_IWL<14884> A_IWL<14883> A_IWL<14882> A_IWL<14881> A_IWL<14880> A_IWL<14879> A_IWL<14878> A_IWL<14877> A_IWL<14876> A_IWL<14875> A_IWL<14874> A_IWL<14873> A_IWL<14872> A_IWL<14871> A_IWL<14870> A_IWL<14869> A_IWL<14868> A_IWL<14867> A_IWL<14866> A_IWL<14865> A_IWL<14864> A_IWL<14863> A_IWL<14862> A_IWL<14861> A_IWL<14860> A_IWL<14859> A_IWL<14858> A_IWL<14857> A_IWL<14856> A_IWL<14855> A_IWL<14854> A_IWL<14853> A_IWL<14852> A_IWL<14851> A_IWL<14850> A_IWL<14849> A_IWL<14848> A_IWL<15871> A_IWL<15870> A_IWL<15869> A_IWL<15868> A_IWL<15867> A_IWL<15866> A_IWL<15865> A_IWL<15864> A_IWL<15863> A_IWL<15862> A_IWL<15861> A_IWL<15860> A_IWL<15859> A_IWL<15858> A_IWL<15857> A_IWL<15856> A_IWL<15855> A_IWL<15854> A_IWL<15853> A_IWL<15852> A_IWL<15851> A_IWL<15850> A_IWL<15849> A_IWL<15848> A_IWL<15847> A_IWL<15846> A_IWL<15845> A_IWL<15844> A_IWL<15843> A_IWL<15842> A_IWL<15841> A_IWL<15840> A_IWL<15839> A_IWL<15838> A_IWL<15837> A_IWL<15836> A_IWL<15835> A_IWL<15834> A_IWL<15833> A_IWL<15832> A_IWL<15831> A_IWL<15830> A_IWL<15829> A_IWL<15828> A_IWL<15827> A_IWL<15826> A_IWL<15825> A_IWL<15824> A_IWL<15823> A_IWL<15822> A_IWL<15821> A_IWL<15820> A_IWL<15819> A_IWL<15818> A_IWL<15817> A_IWL<15816> A_IWL<15815> A_IWL<15814> A_IWL<15813> A_IWL<15812> A_IWL<15811> A_IWL<15810> A_IWL<15809> A_IWL<15808> A_IWL<15807> A_IWL<15806> A_IWL<15805> A_IWL<15804> A_IWL<15803> A_IWL<15802> A_IWL<15801> A_IWL<15800> A_IWL<15799> A_IWL<15798> A_IWL<15797> A_IWL<15796> A_IWL<15795> A_IWL<15794> A_IWL<15793> A_IWL<15792> A_IWL<15791> A_IWL<15790> A_IWL<15789> A_IWL<15788> A_IWL<15787> A_IWL<15786> A_IWL<15785> A_IWL<15784> A_IWL<15783> A_IWL<15782> A_IWL<15781> A_IWL<15780> A_IWL<15779> A_IWL<15778> A_IWL<15777> A_IWL<15776> A_IWL<15775> A_IWL<15774> A_IWL<15773> A_IWL<15772> A_IWL<15771> A_IWL<15770> A_IWL<15769> A_IWL<15768> A_IWL<15767> A_IWL<15766> A_IWL<15765> A_IWL<15764> A_IWL<15763> A_IWL<15762> A_IWL<15761> A_IWL<15760> A_IWL<15759> A_IWL<15758> A_IWL<15757> A_IWL<15756> A_IWL<15755> A_IWL<15754> A_IWL<15753> A_IWL<15752> A_IWL<15751> A_IWL<15750> A_IWL<15749> A_IWL<15748> A_IWL<15747> A_IWL<15746> A_IWL<15745> A_IWL<15744> A_IWL<15743> A_IWL<15742> A_IWL<15741> A_IWL<15740> A_IWL<15739> A_IWL<15738> A_IWL<15737> A_IWL<15736> A_IWL<15735> A_IWL<15734> A_IWL<15733> A_IWL<15732> A_IWL<15731> A_IWL<15730> A_IWL<15729> A_IWL<15728> A_IWL<15727> A_IWL<15726> A_IWL<15725> A_IWL<15724> A_IWL<15723> A_IWL<15722> A_IWL<15721> A_IWL<15720> A_IWL<15719> A_IWL<15718> A_IWL<15717> A_IWL<15716> A_IWL<15715> A_IWL<15714> A_IWL<15713> A_IWL<15712> A_IWL<15711> A_IWL<15710> A_IWL<15709> A_IWL<15708> A_IWL<15707> A_IWL<15706> A_IWL<15705> A_IWL<15704> A_IWL<15703> A_IWL<15702> A_IWL<15701> A_IWL<15700> A_IWL<15699> A_IWL<15698> A_IWL<15697> A_IWL<15696> A_IWL<15695> A_IWL<15694> A_IWL<15693> A_IWL<15692> A_IWL<15691> A_IWL<15690> A_IWL<15689> A_IWL<15688> A_IWL<15687> A_IWL<15686> A_IWL<15685> A_IWL<15684> A_IWL<15683> A_IWL<15682> A_IWL<15681> A_IWL<15680> A_IWL<15679> A_IWL<15678> A_IWL<15677> A_IWL<15676> A_IWL<15675> A_IWL<15674> A_IWL<15673> A_IWL<15672> A_IWL<15671> A_IWL<15670> A_IWL<15669> A_IWL<15668> A_IWL<15667> A_IWL<15666> A_IWL<15665> A_IWL<15664> A_IWL<15663> A_IWL<15662> A_IWL<15661> A_IWL<15660> A_IWL<15659> A_IWL<15658> A_IWL<15657> A_IWL<15656> A_IWL<15655> A_IWL<15654> A_IWL<15653> A_IWL<15652> A_IWL<15651> A_IWL<15650> A_IWL<15649> A_IWL<15648> A_IWL<15647> A_IWL<15646> A_IWL<15645> A_IWL<15644> A_IWL<15643> A_IWL<15642> A_IWL<15641> A_IWL<15640> A_IWL<15639> A_IWL<15638> A_IWL<15637> A_IWL<15636> A_IWL<15635> A_IWL<15634> A_IWL<15633> A_IWL<15632> A_IWL<15631> A_IWL<15630> A_IWL<15629> A_IWL<15628> A_IWL<15627> A_IWL<15626> A_IWL<15625> A_IWL<15624> A_IWL<15623> A_IWL<15622> A_IWL<15621> A_IWL<15620> A_IWL<15619> A_IWL<15618> A_IWL<15617> A_IWL<15616> A_IWL<15615> A_IWL<15614> A_IWL<15613> A_IWL<15612> A_IWL<15611> A_IWL<15610> A_IWL<15609> A_IWL<15608> A_IWL<15607> A_IWL<15606> A_IWL<15605> A_IWL<15604> A_IWL<15603> A_IWL<15602> A_IWL<15601> A_IWL<15600> A_IWL<15599> A_IWL<15598> A_IWL<15597> A_IWL<15596> A_IWL<15595> A_IWL<15594> A_IWL<15593> A_IWL<15592> A_IWL<15591> A_IWL<15590> A_IWL<15589> A_IWL<15588> A_IWL<15587> A_IWL<15586> A_IWL<15585> A_IWL<15584> A_IWL<15583> A_IWL<15582> A_IWL<15581> A_IWL<15580> A_IWL<15579> A_IWL<15578> A_IWL<15577> A_IWL<15576> A_IWL<15575> A_IWL<15574> A_IWL<15573> A_IWL<15572> A_IWL<15571> A_IWL<15570> A_IWL<15569> A_IWL<15568> A_IWL<15567> A_IWL<15566> A_IWL<15565> A_IWL<15564> A_IWL<15563> A_IWL<15562> A_IWL<15561> A_IWL<15560> A_IWL<15559> A_IWL<15558> A_IWL<15557> A_IWL<15556> A_IWL<15555> A_IWL<15554> A_IWL<15553> A_IWL<15552> A_IWL<15551> A_IWL<15550> A_IWL<15549> A_IWL<15548> A_IWL<15547> A_IWL<15546> A_IWL<15545> A_IWL<15544> A_IWL<15543> A_IWL<15542> A_IWL<15541> A_IWL<15540> A_IWL<15539> A_IWL<15538> A_IWL<15537> A_IWL<15536> A_IWL<15535> A_IWL<15534> A_IWL<15533> A_IWL<15532> A_IWL<15531> A_IWL<15530> A_IWL<15529> A_IWL<15528> A_IWL<15527> A_IWL<15526> A_IWL<15525> A_IWL<15524> A_IWL<15523> A_IWL<15522> A_IWL<15521> A_IWL<15520> A_IWL<15519> A_IWL<15518> A_IWL<15517> A_IWL<15516> A_IWL<15515> A_IWL<15514> A_IWL<15513> A_IWL<15512> A_IWL<15511> A_IWL<15510> A_IWL<15509> A_IWL<15508> A_IWL<15507> A_IWL<15506> A_IWL<15505> A_IWL<15504> A_IWL<15503> A_IWL<15502> A_IWL<15501> A_IWL<15500> A_IWL<15499> A_IWL<15498> A_IWL<15497> A_IWL<15496> A_IWL<15495> A_IWL<15494> A_IWL<15493> A_IWL<15492> A_IWL<15491> A_IWL<15490> A_IWL<15489> A_IWL<15488> A_IWL<15487> A_IWL<15486> A_IWL<15485> A_IWL<15484> A_IWL<15483> A_IWL<15482> A_IWL<15481> A_IWL<15480> A_IWL<15479> A_IWL<15478> A_IWL<15477> A_IWL<15476> A_IWL<15475> A_IWL<15474> A_IWL<15473> A_IWL<15472> A_IWL<15471> A_IWL<15470> A_IWL<15469> A_IWL<15468> A_IWL<15467> A_IWL<15466> A_IWL<15465> A_IWL<15464> A_IWL<15463> A_IWL<15462> A_IWL<15461> A_IWL<15460> A_IWL<15459> A_IWL<15458> A_IWL<15457> A_IWL<15456> A_IWL<15455> A_IWL<15454> A_IWL<15453> A_IWL<15452> A_IWL<15451> A_IWL<15450> A_IWL<15449> A_IWL<15448> A_IWL<15447> A_IWL<15446> A_IWL<15445> A_IWL<15444> A_IWL<15443> A_IWL<15442> A_IWL<15441> A_IWL<15440> A_IWL<15439> A_IWL<15438> A_IWL<15437> A_IWL<15436> A_IWL<15435> A_IWL<15434> A_IWL<15433> A_IWL<15432> A_IWL<15431> A_IWL<15430> A_IWL<15429> A_IWL<15428> A_IWL<15427> A_IWL<15426> A_IWL<15425> A_IWL<15424> A_IWL<15423> A_IWL<15422> A_IWL<15421> A_IWL<15420> A_IWL<15419> A_IWL<15418> A_IWL<15417> A_IWL<15416> A_IWL<15415> A_IWL<15414> A_IWL<15413> A_IWL<15412> A_IWL<15411> A_IWL<15410> A_IWL<15409> A_IWL<15408> A_IWL<15407> A_IWL<15406> A_IWL<15405> A_IWL<15404> A_IWL<15403> A_IWL<15402> A_IWL<15401> A_IWL<15400> A_IWL<15399> A_IWL<15398> A_IWL<15397> A_IWL<15396> A_IWL<15395> A_IWL<15394> A_IWL<15393> A_IWL<15392> A_IWL<15391> A_IWL<15390> A_IWL<15389> A_IWL<15388> A_IWL<15387> A_IWL<15386> A_IWL<15385> A_IWL<15384> A_IWL<15383> A_IWL<15382> A_IWL<15381> A_IWL<15380> A_IWL<15379> A_IWL<15378> A_IWL<15377> A_IWL<15376> A_IWL<15375> A_IWL<15374> A_IWL<15373> A_IWL<15372> A_IWL<15371> A_IWL<15370> A_IWL<15369> A_IWL<15368> A_IWL<15367> A_IWL<15366> A_IWL<15365> A_IWL<15364> A_IWL<15363> A_IWL<15362> A_IWL<15361> A_IWL<15360> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<29> A_BLC<59> A_BLC<58> A_BLC_TOP<59> A_BLC_TOP<58> A_BLT<59> A_BLT<58> A_BLT_TOP<59> A_BLT_TOP<58> A_IWL<14847> A_IWL<14846> A_IWL<14845> A_IWL<14844> A_IWL<14843> A_IWL<14842> A_IWL<14841> A_IWL<14840> A_IWL<14839> A_IWL<14838> A_IWL<14837> A_IWL<14836> A_IWL<14835> A_IWL<14834> A_IWL<14833> A_IWL<14832> A_IWL<14831> A_IWL<14830> A_IWL<14829> A_IWL<14828> A_IWL<14827> A_IWL<14826> A_IWL<14825> A_IWL<14824> A_IWL<14823> A_IWL<14822> A_IWL<14821> A_IWL<14820> A_IWL<14819> A_IWL<14818> A_IWL<14817> A_IWL<14816> A_IWL<14815> A_IWL<14814> A_IWL<14813> A_IWL<14812> A_IWL<14811> A_IWL<14810> A_IWL<14809> A_IWL<14808> A_IWL<14807> A_IWL<14806> A_IWL<14805> A_IWL<14804> A_IWL<14803> A_IWL<14802> A_IWL<14801> A_IWL<14800> A_IWL<14799> A_IWL<14798> A_IWL<14797> A_IWL<14796> A_IWL<14795> A_IWL<14794> A_IWL<14793> A_IWL<14792> A_IWL<14791> A_IWL<14790> A_IWL<14789> A_IWL<14788> A_IWL<14787> A_IWL<14786> A_IWL<14785> A_IWL<14784> A_IWL<14783> A_IWL<14782> A_IWL<14781> A_IWL<14780> A_IWL<14779> A_IWL<14778> A_IWL<14777> A_IWL<14776> A_IWL<14775> A_IWL<14774> A_IWL<14773> A_IWL<14772> A_IWL<14771> A_IWL<14770> A_IWL<14769> A_IWL<14768> A_IWL<14767> A_IWL<14766> A_IWL<14765> A_IWL<14764> A_IWL<14763> A_IWL<14762> A_IWL<14761> A_IWL<14760> A_IWL<14759> A_IWL<14758> A_IWL<14757> A_IWL<14756> A_IWL<14755> A_IWL<14754> A_IWL<14753> A_IWL<14752> A_IWL<14751> A_IWL<14750> A_IWL<14749> A_IWL<14748> A_IWL<14747> A_IWL<14746> A_IWL<14745> A_IWL<14744> A_IWL<14743> A_IWL<14742> A_IWL<14741> A_IWL<14740> A_IWL<14739> A_IWL<14738> A_IWL<14737> A_IWL<14736> A_IWL<14735> A_IWL<14734> A_IWL<14733> A_IWL<14732> A_IWL<14731> A_IWL<14730> A_IWL<14729> A_IWL<14728> A_IWL<14727> A_IWL<14726> A_IWL<14725> A_IWL<14724> A_IWL<14723> A_IWL<14722> A_IWL<14721> A_IWL<14720> A_IWL<14719> A_IWL<14718> A_IWL<14717> A_IWL<14716> A_IWL<14715> A_IWL<14714> A_IWL<14713> A_IWL<14712> A_IWL<14711> A_IWL<14710> A_IWL<14709> A_IWL<14708> A_IWL<14707> A_IWL<14706> A_IWL<14705> A_IWL<14704> A_IWL<14703> A_IWL<14702> A_IWL<14701> A_IWL<14700> A_IWL<14699> A_IWL<14698> A_IWL<14697> A_IWL<14696> A_IWL<14695> A_IWL<14694> A_IWL<14693> A_IWL<14692> A_IWL<14691> A_IWL<14690> A_IWL<14689> A_IWL<14688> A_IWL<14687> A_IWL<14686> A_IWL<14685> A_IWL<14684> A_IWL<14683> A_IWL<14682> A_IWL<14681> A_IWL<14680> A_IWL<14679> A_IWL<14678> A_IWL<14677> A_IWL<14676> A_IWL<14675> A_IWL<14674> A_IWL<14673> A_IWL<14672> A_IWL<14671> A_IWL<14670> A_IWL<14669> A_IWL<14668> A_IWL<14667> A_IWL<14666> A_IWL<14665> A_IWL<14664> A_IWL<14663> A_IWL<14662> A_IWL<14661> A_IWL<14660> A_IWL<14659> A_IWL<14658> A_IWL<14657> A_IWL<14656> A_IWL<14655> A_IWL<14654> A_IWL<14653> A_IWL<14652> A_IWL<14651> A_IWL<14650> A_IWL<14649> A_IWL<14648> A_IWL<14647> A_IWL<14646> A_IWL<14645> A_IWL<14644> A_IWL<14643> A_IWL<14642> A_IWL<14641> A_IWL<14640> A_IWL<14639> A_IWL<14638> A_IWL<14637> A_IWL<14636> A_IWL<14635> A_IWL<14634> A_IWL<14633> A_IWL<14632> A_IWL<14631> A_IWL<14630> A_IWL<14629> A_IWL<14628> A_IWL<14627> A_IWL<14626> A_IWL<14625> A_IWL<14624> A_IWL<14623> A_IWL<14622> A_IWL<14621> A_IWL<14620> A_IWL<14619> A_IWL<14618> A_IWL<14617> A_IWL<14616> A_IWL<14615> A_IWL<14614> A_IWL<14613> A_IWL<14612> A_IWL<14611> A_IWL<14610> A_IWL<14609> A_IWL<14608> A_IWL<14607> A_IWL<14606> A_IWL<14605> A_IWL<14604> A_IWL<14603> A_IWL<14602> A_IWL<14601> A_IWL<14600> A_IWL<14599> A_IWL<14598> A_IWL<14597> A_IWL<14596> A_IWL<14595> A_IWL<14594> A_IWL<14593> A_IWL<14592> A_IWL<14591> A_IWL<14590> A_IWL<14589> A_IWL<14588> A_IWL<14587> A_IWL<14586> A_IWL<14585> A_IWL<14584> A_IWL<14583> A_IWL<14582> A_IWL<14581> A_IWL<14580> A_IWL<14579> A_IWL<14578> A_IWL<14577> A_IWL<14576> A_IWL<14575> A_IWL<14574> A_IWL<14573> A_IWL<14572> A_IWL<14571> A_IWL<14570> A_IWL<14569> A_IWL<14568> A_IWL<14567> A_IWL<14566> A_IWL<14565> A_IWL<14564> A_IWL<14563> A_IWL<14562> A_IWL<14561> A_IWL<14560> A_IWL<14559> A_IWL<14558> A_IWL<14557> A_IWL<14556> A_IWL<14555> A_IWL<14554> A_IWL<14553> A_IWL<14552> A_IWL<14551> A_IWL<14550> A_IWL<14549> A_IWL<14548> A_IWL<14547> A_IWL<14546> A_IWL<14545> A_IWL<14544> A_IWL<14543> A_IWL<14542> A_IWL<14541> A_IWL<14540> A_IWL<14539> A_IWL<14538> A_IWL<14537> A_IWL<14536> A_IWL<14535> A_IWL<14534> A_IWL<14533> A_IWL<14532> A_IWL<14531> A_IWL<14530> A_IWL<14529> A_IWL<14528> A_IWL<14527> A_IWL<14526> A_IWL<14525> A_IWL<14524> A_IWL<14523> A_IWL<14522> A_IWL<14521> A_IWL<14520> A_IWL<14519> A_IWL<14518> A_IWL<14517> A_IWL<14516> A_IWL<14515> A_IWL<14514> A_IWL<14513> A_IWL<14512> A_IWL<14511> A_IWL<14510> A_IWL<14509> A_IWL<14508> A_IWL<14507> A_IWL<14506> A_IWL<14505> A_IWL<14504> A_IWL<14503> A_IWL<14502> A_IWL<14501> A_IWL<14500> A_IWL<14499> A_IWL<14498> A_IWL<14497> A_IWL<14496> A_IWL<14495> A_IWL<14494> A_IWL<14493> A_IWL<14492> A_IWL<14491> A_IWL<14490> A_IWL<14489> A_IWL<14488> A_IWL<14487> A_IWL<14486> A_IWL<14485> A_IWL<14484> A_IWL<14483> A_IWL<14482> A_IWL<14481> A_IWL<14480> A_IWL<14479> A_IWL<14478> A_IWL<14477> A_IWL<14476> A_IWL<14475> A_IWL<14474> A_IWL<14473> A_IWL<14472> A_IWL<14471> A_IWL<14470> A_IWL<14469> A_IWL<14468> A_IWL<14467> A_IWL<14466> A_IWL<14465> A_IWL<14464> A_IWL<14463> A_IWL<14462> A_IWL<14461> A_IWL<14460> A_IWL<14459> A_IWL<14458> A_IWL<14457> A_IWL<14456> A_IWL<14455> A_IWL<14454> A_IWL<14453> A_IWL<14452> A_IWL<14451> A_IWL<14450> A_IWL<14449> A_IWL<14448> A_IWL<14447> A_IWL<14446> A_IWL<14445> A_IWL<14444> A_IWL<14443> A_IWL<14442> A_IWL<14441> A_IWL<14440> A_IWL<14439> A_IWL<14438> A_IWL<14437> A_IWL<14436> A_IWL<14435> A_IWL<14434> A_IWL<14433> A_IWL<14432> A_IWL<14431> A_IWL<14430> A_IWL<14429> A_IWL<14428> A_IWL<14427> A_IWL<14426> A_IWL<14425> A_IWL<14424> A_IWL<14423> A_IWL<14422> A_IWL<14421> A_IWL<14420> A_IWL<14419> A_IWL<14418> A_IWL<14417> A_IWL<14416> A_IWL<14415> A_IWL<14414> A_IWL<14413> A_IWL<14412> A_IWL<14411> A_IWL<14410> A_IWL<14409> A_IWL<14408> A_IWL<14407> A_IWL<14406> A_IWL<14405> A_IWL<14404> A_IWL<14403> A_IWL<14402> A_IWL<14401> A_IWL<14400> A_IWL<14399> A_IWL<14398> A_IWL<14397> A_IWL<14396> A_IWL<14395> A_IWL<14394> A_IWL<14393> A_IWL<14392> A_IWL<14391> A_IWL<14390> A_IWL<14389> A_IWL<14388> A_IWL<14387> A_IWL<14386> A_IWL<14385> A_IWL<14384> A_IWL<14383> A_IWL<14382> A_IWL<14381> A_IWL<14380> A_IWL<14379> A_IWL<14378> A_IWL<14377> A_IWL<14376> A_IWL<14375> A_IWL<14374> A_IWL<14373> A_IWL<14372> A_IWL<14371> A_IWL<14370> A_IWL<14369> A_IWL<14368> A_IWL<14367> A_IWL<14366> A_IWL<14365> A_IWL<14364> A_IWL<14363> A_IWL<14362> A_IWL<14361> A_IWL<14360> A_IWL<14359> A_IWL<14358> A_IWL<14357> A_IWL<14356> A_IWL<14355> A_IWL<14354> A_IWL<14353> A_IWL<14352> A_IWL<14351> A_IWL<14350> A_IWL<14349> A_IWL<14348> A_IWL<14347> A_IWL<14346> A_IWL<14345> A_IWL<14344> A_IWL<14343> A_IWL<14342> A_IWL<14341> A_IWL<14340> A_IWL<14339> A_IWL<14338> A_IWL<14337> A_IWL<14336> A_IWL<15359> A_IWL<15358> A_IWL<15357> A_IWL<15356> A_IWL<15355> A_IWL<15354> A_IWL<15353> A_IWL<15352> A_IWL<15351> A_IWL<15350> A_IWL<15349> A_IWL<15348> A_IWL<15347> A_IWL<15346> A_IWL<15345> A_IWL<15344> A_IWL<15343> A_IWL<15342> A_IWL<15341> A_IWL<15340> A_IWL<15339> A_IWL<15338> A_IWL<15337> A_IWL<15336> A_IWL<15335> A_IWL<15334> A_IWL<15333> A_IWL<15332> A_IWL<15331> A_IWL<15330> A_IWL<15329> A_IWL<15328> A_IWL<15327> A_IWL<15326> A_IWL<15325> A_IWL<15324> A_IWL<15323> A_IWL<15322> A_IWL<15321> A_IWL<15320> A_IWL<15319> A_IWL<15318> A_IWL<15317> A_IWL<15316> A_IWL<15315> A_IWL<15314> A_IWL<15313> A_IWL<15312> A_IWL<15311> A_IWL<15310> A_IWL<15309> A_IWL<15308> A_IWL<15307> A_IWL<15306> A_IWL<15305> A_IWL<15304> A_IWL<15303> A_IWL<15302> A_IWL<15301> A_IWL<15300> A_IWL<15299> A_IWL<15298> A_IWL<15297> A_IWL<15296> A_IWL<15295> A_IWL<15294> A_IWL<15293> A_IWL<15292> A_IWL<15291> A_IWL<15290> A_IWL<15289> A_IWL<15288> A_IWL<15287> A_IWL<15286> A_IWL<15285> A_IWL<15284> A_IWL<15283> A_IWL<15282> A_IWL<15281> A_IWL<15280> A_IWL<15279> A_IWL<15278> A_IWL<15277> A_IWL<15276> A_IWL<15275> A_IWL<15274> A_IWL<15273> A_IWL<15272> A_IWL<15271> A_IWL<15270> A_IWL<15269> A_IWL<15268> A_IWL<15267> A_IWL<15266> A_IWL<15265> A_IWL<15264> A_IWL<15263> A_IWL<15262> A_IWL<15261> A_IWL<15260> A_IWL<15259> A_IWL<15258> A_IWL<15257> A_IWL<15256> A_IWL<15255> A_IWL<15254> A_IWL<15253> A_IWL<15252> A_IWL<15251> A_IWL<15250> A_IWL<15249> A_IWL<15248> A_IWL<15247> A_IWL<15246> A_IWL<15245> A_IWL<15244> A_IWL<15243> A_IWL<15242> A_IWL<15241> A_IWL<15240> A_IWL<15239> A_IWL<15238> A_IWL<15237> A_IWL<15236> A_IWL<15235> A_IWL<15234> A_IWL<15233> A_IWL<15232> A_IWL<15231> A_IWL<15230> A_IWL<15229> A_IWL<15228> A_IWL<15227> A_IWL<15226> A_IWL<15225> A_IWL<15224> A_IWL<15223> A_IWL<15222> A_IWL<15221> A_IWL<15220> A_IWL<15219> A_IWL<15218> A_IWL<15217> A_IWL<15216> A_IWL<15215> A_IWL<15214> A_IWL<15213> A_IWL<15212> A_IWL<15211> A_IWL<15210> A_IWL<15209> A_IWL<15208> A_IWL<15207> A_IWL<15206> A_IWL<15205> A_IWL<15204> A_IWL<15203> A_IWL<15202> A_IWL<15201> A_IWL<15200> A_IWL<15199> A_IWL<15198> A_IWL<15197> A_IWL<15196> A_IWL<15195> A_IWL<15194> A_IWL<15193> A_IWL<15192> A_IWL<15191> A_IWL<15190> A_IWL<15189> A_IWL<15188> A_IWL<15187> A_IWL<15186> A_IWL<15185> A_IWL<15184> A_IWL<15183> A_IWL<15182> A_IWL<15181> A_IWL<15180> A_IWL<15179> A_IWL<15178> A_IWL<15177> A_IWL<15176> A_IWL<15175> A_IWL<15174> A_IWL<15173> A_IWL<15172> A_IWL<15171> A_IWL<15170> A_IWL<15169> A_IWL<15168> A_IWL<15167> A_IWL<15166> A_IWL<15165> A_IWL<15164> A_IWL<15163> A_IWL<15162> A_IWL<15161> A_IWL<15160> A_IWL<15159> A_IWL<15158> A_IWL<15157> A_IWL<15156> A_IWL<15155> A_IWL<15154> A_IWL<15153> A_IWL<15152> A_IWL<15151> A_IWL<15150> A_IWL<15149> A_IWL<15148> A_IWL<15147> A_IWL<15146> A_IWL<15145> A_IWL<15144> A_IWL<15143> A_IWL<15142> A_IWL<15141> A_IWL<15140> A_IWL<15139> A_IWL<15138> A_IWL<15137> A_IWL<15136> A_IWL<15135> A_IWL<15134> A_IWL<15133> A_IWL<15132> A_IWL<15131> A_IWL<15130> A_IWL<15129> A_IWL<15128> A_IWL<15127> A_IWL<15126> A_IWL<15125> A_IWL<15124> A_IWL<15123> A_IWL<15122> A_IWL<15121> A_IWL<15120> A_IWL<15119> A_IWL<15118> A_IWL<15117> A_IWL<15116> A_IWL<15115> A_IWL<15114> A_IWL<15113> A_IWL<15112> A_IWL<15111> A_IWL<15110> A_IWL<15109> A_IWL<15108> A_IWL<15107> A_IWL<15106> A_IWL<15105> A_IWL<15104> A_IWL<15103> A_IWL<15102> A_IWL<15101> A_IWL<15100> A_IWL<15099> A_IWL<15098> A_IWL<15097> A_IWL<15096> A_IWL<15095> A_IWL<15094> A_IWL<15093> A_IWL<15092> A_IWL<15091> A_IWL<15090> A_IWL<15089> A_IWL<15088> A_IWL<15087> A_IWL<15086> A_IWL<15085> A_IWL<15084> A_IWL<15083> A_IWL<15082> A_IWL<15081> A_IWL<15080> A_IWL<15079> A_IWL<15078> A_IWL<15077> A_IWL<15076> A_IWL<15075> A_IWL<15074> A_IWL<15073> A_IWL<15072> A_IWL<15071> A_IWL<15070> A_IWL<15069> A_IWL<15068> A_IWL<15067> A_IWL<15066> A_IWL<15065> A_IWL<15064> A_IWL<15063> A_IWL<15062> A_IWL<15061> A_IWL<15060> A_IWL<15059> A_IWL<15058> A_IWL<15057> A_IWL<15056> A_IWL<15055> A_IWL<15054> A_IWL<15053> A_IWL<15052> A_IWL<15051> A_IWL<15050> A_IWL<15049> A_IWL<15048> A_IWL<15047> A_IWL<15046> A_IWL<15045> A_IWL<15044> A_IWL<15043> A_IWL<15042> A_IWL<15041> A_IWL<15040> A_IWL<15039> A_IWL<15038> A_IWL<15037> A_IWL<15036> A_IWL<15035> A_IWL<15034> A_IWL<15033> A_IWL<15032> A_IWL<15031> A_IWL<15030> A_IWL<15029> A_IWL<15028> A_IWL<15027> A_IWL<15026> A_IWL<15025> A_IWL<15024> A_IWL<15023> A_IWL<15022> A_IWL<15021> A_IWL<15020> A_IWL<15019> A_IWL<15018> A_IWL<15017> A_IWL<15016> A_IWL<15015> A_IWL<15014> A_IWL<15013> A_IWL<15012> A_IWL<15011> A_IWL<15010> A_IWL<15009> A_IWL<15008> A_IWL<15007> A_IWL<15006> A_IWL<15005> A_IWL<15004> A_IWL<15003> A_IWL<15002> A_IWL<15001> A_IWL<15000> A_IWL<14999> A_IWL<14998> A_IWL<14997> A_IWL<14996> A_IWL<14995> A_IWL<14994> A_IWL<14993> A_IWL<14992> A_IWL<14991> A_IWL<14990> A_IWL<14989> A_IWL<14988> A_IWL<14987> A_IWL<14986> A_IWL<14985> A_IWL<14984> A_IWL<14983> A_IWL<14982> A_IWL<14981> A_IWL<14980> A_IWL<14979> A_IWL<14978> A_IWL<14977> A_IWL<14976> A_IWL<14975> A_IWL<14974> A_IWL<14973> A_IWL<14972> A_IWL<14971> A_IWL<14970> A_IWL<14969> A_IWL<14968> A_IWL<14967> A_IWL<14966> A_IWL<14965> A_IWL<14964> A_IWL<14963> A_IWL<14962> A_IWL<14961> A_IWL<14960> A_IWL<14959> A_IWL<14958> A_IWL<14957> A_IWL<14956> A_IWL<14955> A_IWL<14954> A_IWL<14953> A_IWL<14952> A_IWL<14951> A_IWL<14950> A_IWL<14949> A_IWL<14948> A_IWL<14947> A_IWL<14946> A_IWL<14945> A_IWL<14944> A_IWL<14943> A_IWL<14942> A_IWL<14941> A_IWL<14940> A_IWL<14939> A_IWL<14938> A_IWL<14937> A_IWL<14936> A_IWL<14935> A_IWL<14934> A_IWL<14933> A_IWL<14932> A_IWL<14931> A_IWL<14930> A_IWL<14929> A_IWL<14928> A_IWL<14927> A_IWL<14926> A_IWL<14925> A_IWL<14924> A_IWL<14923> A_IWL<14922> A_IWL<14921> A_IWL<14920> A_IWL<14919> A_IWL<14918> A_IWL<14917> A_IWL<14916> A_IWL<14915> A_IWL<14914> A_IWL<14913> A_IWL<14912> A_IWL<14911> A_IWL<14910> A_IWL<14909> A_IWL<14908> A_IWL<14907> A_IWL<14906> A_IWL<14905> A_IWL<14904> A_IWL<14903> A_IWL<14902> A_IWL<14901> A_IWL<14900> A_IWL<14899> A_IWL<14898> A_IWL<14897> A_IWL<14896> A_IWL<14895> A_IWL<14894> A_IWL<14893> A_IWL<14892> A_IWL<14891> A_IWL<14890> A_IWL<14889> A_IWL<14888> A_IWL<14887> A_IWL<14886> A_IWL<14885> A_IWL<14884> A_IWL<14883> A_IWL<14882> A_IWL<14881> A_IWL<14880> A_IWL<14879> A_IWL<14878> A_IWL<14877> A_IWL<14876> A_IWL<14875> A_IWL<14874> A_IWL<14873> A_IWL<14872> A_IWL<14871> A_IWL<14870> A_IWL<14869> A_IWL<14868> A_IWL<14867> A_IWL<14866> A_IWL<14865> A_IWL<14864> A_IWL<14863> A_IWL<14862> A_IWL<14861> A_IWL<14860> A_IWL<14859> A_IWL<14858> A_IWL<14857> A_IWL<14856> A_IWL<14855> A_IWL<14854> A_IWL<14853> A_IWL<14852> A_IWL<14851> A_IWL<14850> A_IWL<14849> A_IWL<14848> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<28> A_BLC<57> A_BLC<56> A_BLC_TOP<57> A_BLC_TOP<56> A_BLT<57> A_BLT<56> A_BLT_TOP<57> A_BLT_TOP<56> A_IWL<14335> A_IWL<14334> A_IWL<14333> A_IWL<14332> A_IWL<14331> A_IWL<14330> A_IWL<14329> A_IWL<14328> A_IWL<14327> A_IWL<14326> A_IWL<14325> A_IWL<14324> A_IWL<14323> A_IWL<14322> A_IWL<14321> A_IWL<14320> A_IWL<14319> A_IWL<14318> A_IWL<14317> A_IWL<14316> A_IWL<14315> A_IWL<14314> A_IWL<14313> A_IWL<14312> A_IWL<14311> A_IWL<14310> A_IWL<14309> A_IWL<14308> A_IWL<14307> A_IWL<14306> A_IWL<14305> A_IWL<14304> A_IWL<14303> A_IWL<14302> A_IWL<14301> A_IWL<14300> A_IWL<14299> A_IWL<14298> A_IWL<14297> A_IWL<14296> A_IWL<14295> A_IWL<14294> A_IWL<14293> A_IWL<14292> A_IWL<14291> A_IWL<14290> A_IWL<14289> A_IWL<14288> A_IWL<14287> A_IWL<14286> A_IWL<14285> A_IWL<14284> A_IWL<14283> A_IWL<14282> A_IWL<14281> A_IWL<14280> A_IWL<14279> A_IWL<14278> A_IWL<14277> A_IWL<14276> A_IWL<14275> A_IWL<14274> A_IWL<14273> A_IWL<14272> A_IWL<14271> A_IWL<14270> A_IWL<14269> A_IWL<14268> A_IWL<14267> A_IWL<14266> A_IWL<14265> A_IWL<14264> A_IWL<14263> A_IWL<14262> A_IWL<14261> A_IWL<14260> A_IWL<14259> A_IWL<14258> A_IWL<14257> A_IWL<14256> A_IWL<14255> A_IWL<14254> A_IWL<14253> A_IWL<14252> A_IWL<14251> A_IWL<14250> A_IWL<14249> A_IWL<14248> A_IWL<14247> A_IWL<14246> A_IWL<14245> A_IWL<14244> A_IWL<14243> A_IWL<14242> A_IWL<14241> A_IWL<14240> A_IWL<14239> A_IWL<14238> A_IWL<14237> A_IWL<14236> A_IWL<14235> A_IWL<14234> A_IWL<14233> A_IWL<14232> A_IWL<14231> A_IWL<14230> A_IWL<14229> A_IWL<14228> A_IWL<14227> A_IWL<14226> A_IWL<14225> A_IWL<14224> A_IWL<14223> A_IWL<14222> A_IWL<14221> A_IWL<14220> A_IWL<14219> A_IWL<14218> A_IWL<14217> A_IWL<14216> A_IWL<14215> A_IWL<14214> A_IWL<14213> A_IWL<14212> A_IWL<14211> A_IWL<14210> A_IWL<14209> A_IWL<14208> A_IWL<14207> A_IWL<14206> A_IWL<14205> A_IWL<14204> A_IWL<14203> A_IWL<14202> A_IWL<14201> A_IWL<14200> A_IWL<14199> A_IWL<14198> A_IWL<14197> A_IWL<14196> A_IWL<14195> A_IWL<14194> A_IWL<14193> A_IWL<14192> A_IWL<14191> A_IWL<14190> A_IWL<14189> A_IWL<14188> A_IWL<14187> A_IWL<14186> A_IWL<14185> A_IWL<14184> A_IWL<14183> A_IWL<14182> A_IWL<14181> A_IWL<14180> A_IWL<14179> A_IWL<14178> A_IWL<14177> A_IWL<14176> A_IWL<14175> A_IWL<14174> A_IWL<14173> A_IWL<14172> A_IWL<14171> A_IWL<14170> A_IWL<14169> A_IWL<14168> A_IWL<14167> A_IWL<14166> A_IWL<14165> A_IWL<14164> A_IWL<14163> A_IWL<14162> A_IWL<14161> A_IWL<14160> A_IWL<14159> A_IWL<14158> A_IWL<14157> A_IWL<14156> A_IWL<14155> A_IWL<14154> A_IWL<14153> A_IWL<14152> A_IWL<14151> A_IWL<14150> A_IWL<14149> A_IWL<14148> A_IWL<14147> A_IWL<14146> A_IWL<14145> A_IWL<14144> A_IWL<14143> A_IWL<14142> A_IWL<14141> A_IWL<14140> A_IWL<14139> A_IWL<14138> A_IWL<14137> A_IWL<14136> A_IWL<14135> A_IWL<14134> A_IWL<14133> A_IWL<14132> A_IWL<14131> A_IWL<14130> A_IWL<14129> A_IWL<14128> A_IWL<14127> A_IWL<14126> A_IWL<14125> A_IWL<14124> A_IWL<14123> A_IWL<14122> A_IWL<14121> A_IWL<14120> A_IWL<14119> A_IWL<14118> A_IWL<14117> A_IWL<14116> A_IWL<14115> A_IWL<14114> A_IWL<14113> A_IWL<14112> A_IWL<14111> A_IWL<14110> A_IWL<14109> A_IWL<14108> A_IWL<14107> A_IWL<14106> A_IWL<14105> A_IWL<14104> A_IWL<14103> A_IWL<14102> A_IWL<14101> A_IWL<14100> A_IWL<14099> A_IWL<14098> A_IWL<14097> A_IWL<14096> A_IWL<14095> A_IWL<14094> A_IWL<14093> A_IWL<14092> A_IWL<14091> A_IWL<14090> A_IWL<14089> A_IWL<14088> A_IWL<14087> A_IWL<14086> A_IWL<14085> A_IWL<14084> A_IWL<14083> A_IWL<14082> A_IWL<14081> A_IWL<14080> A_IWL<14079> A_IWL<14078> A_IWL<14077> A_IWL<14076> A_IWL<14075> A_IWL<14074> A_IWL<14073> A_IWL<14072> A_IWL<14071> A_IWL<14070> A_IWL<14069> A_IWL<14068> A_IWL<14067> A_IWL<14066> A_IWL<14065> A_IWL<14064> A_IWL<14063> A_IWL<14062> A_IWL<14061> A_IWL<14060> A_IWL<14059> A_IWL<14058> A_IWL<14057> A_IWL<14056> A_IWL<14055> A_IWL<14054> A_IWL<14053> A_IWL<14052> A_IWL<14051> A_IWL<14050> A_IWL<14049> A_IWL<14048> A_IWL<14047> A_IWL<14046> A_IWL<14045> A_IWL<14044> A_IWL<14043> A_IWL<14042> A_IWL<14041> A_IWL<14040> A_IWL<14039> A_IWL<14038> A_IWL<14037> A_IWL<14036> A_IWL<14035> A_IWL<14034> A_IWL<14033> A_IWL<14032> A_IWL<14031> A_IWL<14030> A_IWL<14029> A_IWL<14028> A_IWL<14027> A_IWL<14026> A_IWL<14025> A_IWL<14024> A_IWL<14023> A_IWL<14022> A_IWL<14021> A_IWL<14020> A_IWL<14019> A_IWL<14018> A_IWL<14017> A_IWL<14016> A_IWL<14015> A_IWL<14014> A_IWL<14013> A_IWL<14012> A_IWL<14011> A_IWL<14010> A_IWL<14009> A_IWL<14008> A_IWL<14007> A_IWL<14006> A_IWL<14005> A_IWL<14004> A_IWL<14003> A_IWL<14002> A_IWL<14001> A_IWL<14000> A_IWL<13999> A_IWL<13998> A_IWL<13997> A_IWL<13996> A_IWL<13995> A_IWL<13994> A_IWL<13993> A_IWL<13992> A_IWL<13991> A_IWL<13990> A_IWL<13989> A_IWL<13988> A_IWL<13987> A_IWL<13986> A_IWL<13985> A_IWL<13984> A_IWL<13983> A_IWL<13982> A_IWL<13981> A_IWL<13980> A_IWL<13979> A_IWL<13978> A_IWL<13977> A_IWL<13976> A_IWL<13975> A_IWL<13974> A_IWL<13973> A_IWL<13972> A_IWL<13971> A_IWL<13970> A_IWL<13969> A_IWL<13968> A_IWL<13967> A_IWL<13966> A_IWL<13965> A_IWL<13964> A_IWL<13963> A_IWL<13962> A_IWL<13961> A_IWL<13960> A_IWL<13959> A_IWL<13958> A_IWL<13957> A_IWL<13956> A_IWL<13955> A_IWL<13954> A_IWL<13953> A_IWL<13952> A_IWL<13951> A_IWL<13950> A_IWL<13949> A_IWL<13948> A_IWL<13947> A_IWL<13946> A_IWL<13945> A_IWL<13944> A_IWL<13943> A_IWL<13942> A_IWL<13941> A_IWL<13940> A_IWL<13939> A_IWL<13938> A_IWL<13937> A_IWL<13936> A_IWL<13935> A_IWL<13934> A_IWL<13933> A_IWL<13932> A_IWL<13931> A_IWL<13930> A_IWL<13929> A_IWL<13928> A_IWL<13927> A_IWL<13926> A_IWL<13925> A_IWL<13924> A_IWL<13923> A_IWL<13922> A_IWL<13921> A_IWL<13920> A_IWL<13919> A_IWL<13918> A_IWL<13917> A_IWL<13916> A_IWL<13915> A_IWL<13914> A_IWL<13913> A_IWL<13912> A_IWL<13911> A_IWL<13910> A_IWL<13909> A_IWL<13908> A_IWL<13907> A_IWL<13906> A_IWL<13905> A_IWL<13904> A_IWL<13903> A_IWL<13902> A_IWL<13901> A_IWL<13900> A_IWL<13899> A_IWL<13898> A_IWL<13897> A_IWL<13896> A_IWL<13895> A_IWL<13894> A_IWL<13893> A_IWL<13892> A_IWL<13891> A_IWL<13890> A_IWL<13889> A_IWL<13888> A_IWL<13887> A_IWL<13886> A_IWL<13885> A_IWL<13884> A_IWL<13883> A_IWL<13882> A_IWL<13881> A_IWL<13880> A_IWL<13879> A_IWL<13878> A_IWL<13877> A_IWL<13876> A_IWL<13875> A_IWL<13874> A_IWL<13873> A_IWL<13872> A_IWL<13871> A_IWL<13870> A_IWL<13869> A_IWL<13868> A_IWL<13867> A_IWL<13866> A_IWL<13865> A_IWL<13864> A_IWL<13863> A_IWL<13862> A_IWL<13861> A_IWL<13860> A_IWL<13859> A_IWL<13858> A_IWL<13857> A_IWL<13856> A_IWL<13855> A_IWL<13854> A_IWL<13853> A_IWL<13852> A_IWL<13851> A_IWL<13850> A_IWL<13849> A_IWL<13848> A_IWL<13847> A_IWL<13846> A_IWL<13845> A_IWL<13844> A_IWL<13843> A_IWL<13842> A_IWL<13841> A_IWL<13840> A_IWL<13839> A_IWL<13838> A_IWL<13837> A_IWL<13836> A_IWL<13835> A_IWL<13834> A_IWL<13833> A_IWL<13832> A_IWL<13831> A_IWL<13830> A_IWL<13829> A_IWL<13828> A_IWL<13827> A_IWL<13826> A_IWL<13825> A_IWL<13824> A_IWL<14847> A_IWL<14846> A_IWL<14845> A_IWL<14844> A_IWL<14843> A_IWL<14842> A_IWL<14841> A_IWL<14840> A_IWL<14839> A_IWL<14838> A_IWL<14837> A_IWL<14836> A_IWL<14835> A_IWL<14834> A_IWL<14833> A_IWL<14832> A_IWL<14831> A_IWL<14830> A_IWL<14829> A_IWL<14828> A_IWL<14827> A_IWL<14826> A_IWL<14825> A_IWL<14824> A_IWL<14823> A_IWL<14822> A_IWL<14821> A_IWL<14820> A_IWL<14819> A_IWL<14818> A_IWL<14817> A_IWL<14816> A_IWL<14815> A_IWL<14814> A_IWL<14813> A_IWL<14812> A_IWL<14811> A_IWL<14810> A_IWL<14809> A_IWL<14808> A_IWL<14807> A_IWL<14806> A_IWL<14805> A_IWL<14804> A_IWL<14803> A_IWL<14802> A_IWL<14801> A_IWL<14800> A_IWL<14799> A_IWL<14798> A_IWL<14797> A_IWL<14796> A_IWL<14795> A_IWL<14794> A_IWL<14793> A_IWL<14792> A_IWL<14791> A_IWL<14790> A_IWL<14789> A_IWL<14788> A_IWL<14787> A_IWL<14786> A_IWL<14785> A_IWL<14784> A_IWL<14783> A_IWL<14782> A_IWL<14781> A_IWL<14780> A_IWL<14779> A_IWL<14778> A_IWL<14777> A_IWL<14776> A_IWL<14775> A_IWL<14774> A_IWL<14773> A_IWL<14772> A_IWL<14771> A_IWL<14770> A_IWL<14769> A_IWL<14768> A_IWL<14767> A_IWL<14766> A_IWL<14765> A_IWL<14764> A_IWL<14763> A_IWL<14762> A_IWL<14761> A_IWL<14760> A_IWL<14759> A_IWL<14758> A_IWL<14757> A_IWL<14756> A_IWL<14755> A_IWL<14754> A_IWL<14753> A_IWL<14752> A_IWL<14751> A_IWL<14750> A_IWL<14749> A_IWL<14748> A_IWL<14747> A_IWL<14746> A_IWL<14745> A_IWL<14744> A_IWL<14743> A_IWL<14742> A_IWL<14741> A_IWL<14740> A_IWL<14739> A_IWL<14738> A_IWL<14737> A_IWL<14736> A_IWL<14735> A_IWL<14734> A_IWL<14733> A_IWL<14732> A_IWL<14731> A_IWL<14730> A_IWL<14729> A_IWL<14728> A_IWL<14727> A_IWL<14726> A_IWL<14725> A_IWL<14724> A_IWL<14723> A_IWL<14722> A_IWL<14721> A_IWL<14720> A_IWL<14719> A_IWL<14718> A_IWL<14717> A_IWL<14716> A_IWL<14715> A_IWL<14714> A_IWL<14713> A_IWL<14712> A_IWL<14711> A_IWL<14710> A_IWL<14709> A_IWL<14708> A_IWL<14707> A_IWL<14706> A_IWL<14705> A_IWL<14704> A_IWL<14703> A_IWL<14702> A_IWL<14701> A_IWL<14700> A_IWL<14699> A_IWL<14698> A_IWL<14697> A_IWL<14696> A_IWL<14695> A_IWL<14694> A_IWL<14693> A_IWL<14692> A_IWL<14691> A_IWL<14690> A_IWL<14689> A_IWL<14688> A_IWL<14687> A_IWL<14686> A_IWL<14685> A_IWL<14684> A_IWL<14683> A_IWL<14682> A_IWL<14681> A_IWL<14680> A_IWL<14679> A_IWL<14678> A_IWL<14677> A_IWL<14676> A_IWL<14675> A_IWL<14674> A_IWL<14673> A_IWL<14672> A_IWL<14671> A_IWL<14670> A_IWL<14669> A_IWL<14668> A_IWL<14667> A_IWL<14666> A_IWL<14665> A_IWL<14664> A_IWL<14663> A_IWL<14662> A_IWL<14661> A_IWL<14660> A_IWL<14659> A_IWL<14658> A_IWL<14657> A_IWL<14656> A_IWL<14655> A_IWL<14654> A_IWL<14653> A_IWL<14652> A_IWL<14651> A_IWL<14650> A_IWL<14649> A_IWL<14648> A_IWL<14647> A_IWL<14646> A_IWL<14645> A_IWL<14644> A_IWL<14643> A_IWL<14642> A_IWL<14641> A_IWL<14640> A_IWL<14639> A_IWL<14638> A_IWL<14637> A_IWL<14636> A_IWL<14635> A_IWL<14634> A_IWL<14633> A_IWL<14632> A_IWL<14631> A_IWL<14630> A_IWL<14629> A_IWL<14628> A_IWL<14627> A_IWL<14626> A_IWL<14625> A_IWL<14624> A_IWL<14623> A_IWL<14622> A_IWL<14621> A_IWL<14620> A_IWL<14619> A_IWL<14618> A_IWL<14617> A_IWL<14616> A_IWL<14615> A_IWL<14614> A_IWL<14613> A_IWL<14612> A_IWL<14611> A_IWL<14610> A_IWL<14609> A_IWL<14608> A_IWL<14607> A_IWL<14606> A_IWL<14605> A_IWL<14604> A_IWL<14603> A_IWL<14602> A_IWL<14601> A_IWL<14600> A_IWL<14599> A_IWL<14598> A_IWL<14597> A_IWL<14596> A_IWL<14595> A_IWL<14594> A_IWL<14593> A_IWL<14592> A_IWL<14591> A_IWL<14590> A_IWL<14589> A_IWL<14588> A_IWL<14587> A_IWL<14586> A_IWL<14585> A_IWL<14584> A_IWL<14583> A_IWL<14582> A_IWL<14581> A_IWL<14580> A_IWL<14579> A_IWL<14578> A_IWL<14577> A_IWL<14576> A_IWL<14575> A_IWL<14574> A_IWL<14573> A_IWL<14572> A_IWL<14571> A_IWL<14570> A_IWL<14569> A_IWL<14568> A_IWL<14567> A_IWL<14566> A_IWL<14565> A_IWL<14564> A_IWL<14563> A_IWL<14562> A_IWL<14561> A_IWL<14560> A_IWL<14559> A_IWL<14558> A_IWL<14557> A_IWL<14556> A_IWL<14555> A_IWL<14554> A_IWL<14553> A_IWL<14552> A_IWL<14551> A_IWL<14550> A_IWL<14549> A_IWL<14548> A_IWL<14547> A_IWL<14546> A_IWL<14545> A_IWL<14544> A_IWL<14543> A_IWL<14542> A_IWL<14541> A_IWL<14540> A_IWL<14539> A_IWL<14538> A_IWL<14537> A_IWL<14536> A_IWL<14535> A_IWL<14534> A_IWL<14533> A_IWL<14532> A_IWL<14531> A_IWL<14530> A_IWL<14529> A_IWL<14528> A_IWL<14527> A_IWL<14526> A_IWL<14525> A_IWL<14524> A_IWL<14523> A_IWL<14522> A_IWL<14521> A_IWL<14520> A_IWL<14519> A_IWL<14518> A_IWL<14517> A_IWL<14516> A_IWL<14515> A_IWL<14514> A_IWL<14513> A_IWL<14512> A_IWL<14511> A_IWL<14510> A_IWL<14509> A_IWL<14508> A_IWL<14507> A_IWL<14506> A_IWL<14505> A_IWL<14504> A_IWL<14503> A_IWL<14502> A_IWL<14501> A_IWL<14500> A_IWL<14499> A_IWL<14498> A_IWL<14497> A_IWL<14496> A_IWL<14495> A_IWL<14494> A_IWL<14493> A_IWL<14492> A_IWL<14491> A_IWL<14490> A_IWL<14489> A_IWL<14488> A_IWL<14487> A_IWL<14486> A_IWL<14485> A_IWL<14484> A_IWL<14483> A_IWL<14482> A_IWL<14481> A_IWL<14480> A_IWL<14479> A_IWL<14478> A_IWL<14477> A_IWL<14476> A_IWL<14475> A_IWL<14474> A_IWL<14473> A_IWL<14472> A_IWL<14471> A_IWL<14470> A_IWL<14469> A_IWL<14468> A_IWL<14467> A_IWL<14466> A_IWL<14465> A_IWL<14464> A_IWL<14463> A_IWL<14462> A_IWL<14461> A_IWL<14460> A_IWL<14459> A_IWL<14458> A_IWL<14457> A_IWL<14456> A_IWL<14455> A_IWL<14454> A_IWL<14453> A_IWL<14452> A_IWL<14451> A_IWL<14450> A_IWL<14449> A_IWL<14448> A_IWL<14447> A_IWL<14446> A_IWL<14445> A_IWL<14444> A_IWL<14443> A_IWL<14442> A_IWL<14441> A_IWL<14440> A_IWL<14439> A_IWL<14438> A_IWL<14437> A_IWL<14436> A_IWL<14435> A_IWL<14434> A_IWL<14433> A_IWL<14432> A_IWL<14431> A_IWL<14430> A_IWL<14429> A_IWL<14428> A_IWL<14427> A_IWL<14426> A_IWL<14425> A_IWL<14424> A_IWL<14423> A_IWL<14422> A_IWL<14421> A_IWL<14420> A_IWL<14419> A_IWL<14418> A_IWL<14417> A_IWL<14416> A_IWL<14415> A_IWL<14414> A_IWL<14413> A_IWL<14412> A_IWL<14411> A_IWL<14410> A_IWL<14409> A_IWL<14408> A_IWL<14407> A_IWL<14406> A_IWL<14405> A_IWL<14404> A_IWL<14403> A_IWL<14402> A_IWL<14401> A_IWL<14400> A_IWL<14399> A_IWL<14398> A_IWL<14397> A_IWL<14396> A_IWL<14395> A_IWL<14394> A_IWL<14393> A_IWL<14392> A_IWL<14391> A_IWL<14390> A_IWL<14389> A_IWL<14388> A_IWL<14387> A_IWL<14386> A_IWL<14385> A_IWL<14384> A_IWL<14383> A_IWL<14382> A_IWL<14381> A_IWL<14380> A_IWL<14379> A_IWL<14378> A_IWL<14377> A_IWL<14376> A_IWL<14375> A_IWL<14374> A_IWL<14373> A_IWL<14372> A_IWL<14371> A_IWL<14370> A_IWL<14369> A_IWL<14368> A_IWL<14367> A_IWL<14366> A_IWL<14365> A_IWL<14364> A_IWL<14363> A_IWL<14362> A_IWL<14361> A_IWL<14360> A_IWL<14359> A_IWL<14358> A_IWL<14357> A_IWL<14356> A_IWL<14355> A_IWL<14354> A_IWL<14353> A_IWL<14352> A_IWL<14351> A_IWL<14350> A_IWL<14349> A_IWL<14348> A_IWL<14347> A_IWL<14346> A_IWL<14345> A_IWL<14344> A_IWL<14343> A_IWL<14342> A_IWL<14341> A_IWL<14340> A_IWL<14339> A_IWL<14338> A_IWL<14337> A_IWL<14336> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<27> A_BLC<55> A_BLC<54> A_BLC_TOP<55> A_BLC_TOP<54> A_BLT<55> A_BLT<54> A_BLT_TOP<55> A_BLT_TOP<54> A_IWL<13823> A_IWL<13822> A_IWL<13821> A_IWL<13820> A_IWL<13819> A_IWL<13818> A_IWL<13817> A_IWL<13816> A_IWL<13815> A_IWL<13814> A_IWL<13813> A_IWL<13812> A_IWL<13811> A_IWL<13810> A_IWL<13809> A_IWL<13808> A_IWL<13807> A_IWL<13806> A_IWL<13805> A_IWL<13804> A_IWL<13803> A_IWL<13802> A_IWL<13801> A_IWL<13800> A_IWL<13799> A_IWL<13798> A_IWL<13797> A_IWL<13796> A_IWL<13795> A_IWL<13794> A_IWL<13793> A_IWL<13792> A_IWL<13791> A_IWL<13790> A_IWL<13789> A_IWL<13788> A_IWL<13787> A_IWL<13786> A_IWL<13785> A_IWL<13784> A_IWL<13783> A_IWL<13782> A_IWL<13781> A_IWL<13780> A_IWL<13779> A_IWL<13778> A_IWL<13777> A_IWL<13776> A_IWL<13775> A_IWL<13774> A_IWL<13773> A_IWL<13772> A_IWL<13771> A_IWL<13770> A_IWL<13769> A_IWL<13768> A_IWL<13767> A_IWL<13766> A_IWL<13765> A_IWL<13764> A_IWL<13763> A_IWL<13762> A_IWL<13761> A_IWL<13760> A_IWL<13759> A_IWL<13758> A_IWL<13757> A_IWL<13756> A_IWL<13755> A_IWL<13754> A_IWL<13753> A_IWL<13752> A_IWL<13751> A_IWL<13750> A_IWL<13749> A_IWL<13748> A_IWL<13747> A_IWL<13746> A_IWL<13745> A_IWL<13744> A_IWL<13743> A_IWL<13742> A_IWL<13741> A_IWL<13740> A_IWL<13739> A_IWL<13738> A_IWL<13737> A_IWL<13736> A_IWL<13735> A_IWL<13734> A_IWL<13733> A_IWL<13732> A_IWL<13731> A_IWL<13730> A_IWL<13729> A_IWL<13728> A_IWL<13727> A_IWL<13726> A_IWL<13725> A_IWL<13724> A_IWL<13723> A_IWL<13722> A_IWL<13721> A_IWL<13720> A_IWL<13719> A_IWL<13718> A_IWL<13717> A_IWL<13716> A_IWL<13715> A_IWL<13714> A_IWL<13713> A_IWL<13712> A_IWL<13711> A_IWL<13710> A_IWL<13709> A_IWL<13708> A_IWL<13707> A_IWL<13706> A_IWL<13705> A_IWL<13704> A_IWL<13703> A_IWL<13702> A_IWL<13701> A_IWL<13700> A_IWL<13699> A_IWL<13698> A_IWL<13697> A_IWL<13696> A_IWL<13695> A_IWL<13694> A_IWL<13693> A_IWL<13692> A_IWL<13691> A_IWL<13690> A_IWL<13689> A_IWL<13688> A_IWL<13687> A_IWL<13686> A_IWL<13685> A_IWL<13684> A_IWL<13683> A_IWL<13682> A_IWL<13681> A_IWL<13680> A_IWL<13679> A_IWL<13678> A_IWL<13677> A_IWL<13676> A_IWL<13675> A_IWL<13674> A_IWL<13673> A_IWL<13672> A_IWL<13671> A_IWL<13670> A_IWL<13669> A_IWL<13668> A_IWL<13667> A_IWL<13666> A_IWL<13665> A_IWL<13664> A_IWL<13663> A_IWL<13662> A_IWL<13661> A_IWL<13660> A_IWL<13659> A_IWL<13658> A_IWL<13657> A_IWL<13656> A_IWL<13655> A_IWL<13654> A_IWL<13653> A_IWL<13652> A_IWL<13651> A_IWL<13650> A_IWL<13649> A_IWL<13648> A_IWL<13647> A_IWL<13646> A_IWL<13645> A_IWL<13644> A_IWL<13643> A_IWL<13642> A_IWL<13641> A_IWL<13640> A_IWL<13639> A_IWL<13638> A_IWL<13637> A_IWL<13636> A_IWL<13635> A_IWL<13634> A_IWL<13633> A_IWL<13632> A_IWL<13631> A_IWL<13630> A_IWL<13629> A_IWL<13628> A_IWL<13627> A_IWL<13626> A_IWL<13625> A_IWL<13624> A_IWL<13623> A_IWL<13622> A_IWL<13621> A_IWL<13620> A_IWL<13619> A_IWL<13618> A_IWL<13617> A_IWL<13616> A_IWL<13615> A_IWL<13614> A_IWL<13613> A_IWL<13612> A_IWL<13611> A_IWL<13610> A_IWL<13609> A_IWL<13608> A_IWL<13607> A_IWL<13606> A_IWL<13605> A_IWL<13604> A_IWL<13603> A_IWL<13602> A_IWL<13601> A_IWL<13600> A_IWL<13599> A_IWL<13598> A_IWL<13597> A_IWL<13596> A_IWL<13595> A_IWL<13594> A_IWL<13593> A_IWL<13592> A_IWL<13591> A_IWL<13590> A_IWL<13589> A_IWL<13588> A_IWL<13587> A_IWL<13586> A_IWL<13585> A_IWL<13584> A_IWL<13583> A_IWL<13582> A_IWL<13581> A_IWL<13580> A_IWL<13579> A_IWL<13578> A_IWL<13577> A_IWL<13576> A_IWL<13575> A_IWL<13574> A_IWL<13573> A_IWL<13572> A_IWL<13571> A_IWL<13570> A_IWL<13569> A_IWL<13568> A_IWL<13567> A_IWL<13566> A_IWL<13565> A_IWL<13564> A_IWL<13563> A_IWL<13562> A_IWL<13561> A_IWL<13560> A_IWL<13559> A_IWL<13558> A_IWL<13557> A_IWL<13556> A_IWL<13555> A_IWL<13554> A_IWL<13553> A_IWL<13552> A_IWL<13551> A_IWL<13550> A_IWL<13549> A_IWL<13548> A_IWL<13547> A_IWL<13546> A_IWL<13545> A_IWL<13544> A_IWL<13543> A_IWL<13542> A_IWL<13541> A_IWL<13540> A_IWL<13539> A_IWL<13538> A_IWL<13537> A_IWL<13536> A_IWL<13535> A_IWL<13534> A_IWL<13533> A_IWL<13532> A_IWL<13531> A_IWL<13530> A_IWL<13529> A_IWL<13528> A_IWL<13527> A_IWL<13526> A_IWL<13525> A_IWL<13524> A_IWL<13523> A_IWL<13522> A_IWL<13521> A_IWL<13520> A_IWL<13519> A_IWL<13518> A_IWL<13517> A_IWL<13516> A_IWL<13515> A_IWL<13514> A_IWL<13513> A_IWL<13512> A_IWL<13511> A_IWL<13510> A_IWL<13509> A_IWL<13508> A_IWL<13507> A_IWL<13506> A_IWL<13505> A_IWL<13504> A_IWL<13503> A_IWL<13502> A_IWL<13501> A_IWL<13500> A_IWL<13499> A_IWL<13498> A_IWL<13497> A_IWL<13496> A_IWL<13495> A_IWL<13494> A_IWL<13493> A_IWL<13492> A_IWL<13491> A_IWL<13490> A_IWL<13489> A_IWL<13488> A_IWL<13487> A_IWL<13486> A_IWL<13485> A_IWL<13484> A_IWL<13483> A_IWL<13482> A_IWL<13481> A_IWL<13480> A_IWL<13479> A_IWL<13478> A_IWL<13477> A_IWL<13476> A_IWL<13475> A_IWL<13474> A_IWL<13473> A_IWL<13472> A_IWL<13471> A_IWL<13470> A_IWL<13469> A_IWL<13468> A_IWL<13467> A_IWL<13466> A_IWL<13465> A_IWL<13464> A_IWL<13463> A_IWL<13462> A_IWL<13461> A_IWL<13460> A_IWL<13459> A_IWL<13458> A_IWL<13457> A_IWL<13456> A_IWL<13455> A_IWL<13454> A_IWL<13453> A_IWL<13452> A_IWL<13451> A_IWL<13450> A_IWL<13449> A_IWL<13448> A_IWL<13447> A_IWL<13446> A_IWL<13445> A_IWL<13444> A_IWL<13443> A_IWL<13442> A_IWL<13441> A_IWL<13440> A_IWL<13439> A_IWL<13438> A_IWL<13437> A_IWL<13436> A_IWL<13435> A_IWL<13434> A_IWL<13433> A_IWL<13432> A_IWL<13431> A_IWL<13430> A_IWL<13429> A_IWL<13428> A_IWL<13427> A_IWL<13426> A_IWL<13425> A_IWL<13424> A_IWL<13423> A_IWL<13422> A_IWL<13421> A_IWL<13420> A_IWL<13419> A_IWL<13418> A_IWL<13417> A_IWL<13416> A_IWL<13415> A_IWL<13414> A_IWL<13413> A_IWL<13412> A_IWL<13411> A_IWL<13410> A_IWL<13409> A_IWL<13408> A_IWL<13407> A_IWL<13406> A_IWL<13405> A_IWL<13404> A_IWL<13403> A_IWL<13402> A_IWL<13401> A_IWL<13400> A_IWL<13399> A_IWL<13398> A_IWL<13397> A_IWL<13396> A_IWL<13395> A_IWL<13394> A_IWL<13393> A_IWL<13392> A_IWL<13391> A_IWL<13390> A_IWL<13389> A_IWL<13388> A_IWL<13387> A_IWL<13386> A_IWL<13385> A_IWL<13384> A_IWL<13383> A_IWL<13382> A_IWL<13381> A_IWL<13380> A_IWL<13379> A_IWL<13378> A_IWL<13377> A_IWL<13376> A_IWL<13375> A_IWL<13374> A_IWL<13373> A_IWL<13372> A_IWL<13371> A_IWL<13370> A_IWL<13369> A_IWL<13368> A_IWL<13367> A_IWL<13366> A_IWL<13365> A_IWL<13364> A_IWL<13363> A_IWL<13362> A_IWL<13361> A_IWL<13360> A_IWL<13359> A_IWL<13358> A_IWL<13357> A_IWL<13356> A_IWL<13355> A_IWL<13354> A_IWL<13353> A_IWL<13352> A_IWL<13351> A_IWL<13350> A_IWL<13349> A_IWL<13348> A_IWL<13347> A_IWL<13346> A_IWL<13345> A_IWL<13344> A_IWL<13343> A_IWL<13342> A_IWL<13341> A_IWL<13340> A_IWL<13339> A_IWL<13338> A_IWL<13337> A_IWL<13336> A_IWL<13335> A_IWL<13334> A_IWL<13333> A_IWL<13332> A_IWL<13331> A_IWL<13330> A_IWL<13329> A_IWL<13328> A_IWL<13327> A_IWL<13326> A_IWL<13325> A_IWL<13324> A_IWL<13323> A_IWL<13322> A_IWL<13321> A_IWL<13320> A_IWL<13319> A_IWL<13318> A_IWL<13317> A_IWL<13316> A_IWL<13315> A_IWL<13314> A_IWL<13313> A_IWL<13312> A_IWL<14335> A_IWL<14334> A_IWL<14333> A_IWL<14332> A_IWL<14331> A_IWL<14330> A_IWL<14329> A_IWL<14328> A_IWL<14327> A_IWL<14326> A_IWL<14325> A_IWL<14324> A_IWL<14323> A_IWL<14322> A_IWL<14321> A_IWL<14320> A_IWL<14319> A_IWL<14318> A_IWL<14317> A_IWL<14316> A_IWL<14315> A_IWL<14314> A_IWL<14313> A_IWL<14312> A_IWL<14311> A_IWL<14310> A_IWL<14309> A_IWL<14308> A_IWL<14307> A_IWL<14306> A_IWL<14305> A_IWL<14304> A_IWL<14303> A_IWL<14302> A_IWL<14301> A_IWL<14300> A_IWL<14299> A_IWL<14298> A_IWL<14297> A_IWL<14296> A_IWL<14295> A_IWL<14294> A_IWL<14293> A_IWL<14292> A_IWL<14291> A_IWL<14290> A_IWL<14289> A_IWL<14288> A_IWL<14287> A_IWL<14286> A_IWL<14285> A_IWL<14284> A_IWL<14283> A_IWL<14282> A_IWL<14281> A_IWL<14280> A_IWL<14279> A_IWL<14278> A_IWL<14277> A_IWL<14276> A_IWL<14275> A_IWL<14274> A_IWL<14273> A_IWL<14272> A_IWL<14271> A_IWL<14270> A_IWL<14269> A_IWL<14268> A_IWL<14267> A_IWL<14266> A_IWL<14265> A_IWL<14264> A_IWL<14263> A_IWL<14262> A_IWL<14261> A_IWL<14260> A_IWL<14259> A_IWL<14258> A_IWL<14257> A_IWL<14256> A_IWL<14255> A_IWL<14254> A_IWL<14253> A_IWL<14252> A_IWL<14251> A_IWL<14250> A_IWL<14249> A_IWL<14248> A_IWL<14247> A_IWL<14246> A_IWL<14245> A_IWL<14244> A_IWL<14243> A_IWL<14242> A_IWL<14241> A_IWL<14240> A_IWL<14239> A_IWL<14238> A_IWL<14237> A_IWL<14236> A_IWL<14235> A_IWL<14234> A_IWL<14233> A_IWL<14232> A_IWL<14231> A_IWL<14230> A_IWL<14229> A_IWL<14228> A_IWL<14227> A_IWL<14226> A_IWL<14225> A_IWL<14224> A_IWL<14223> A_IWL<14222> A_IWL<14221> A_IWL<14220> A_IWL<14219> A_IWL<14218> A_IWL<14217> A_IWL<14216> A_IWL<14215> A_IWL<14214> A_IWL<14213> A_IWL<14212> A_IWL<14211> A_IWL<14210> A_IWL<14209> A_IWL<14208> A_IWL<14207> A_IWL<14206> A_IWL<14205> A_IWL<14204> A_IWL<14203> A_IWL<14202> A_IWL<14201> A_IWL<14200> A_IWL<14199> A_IWL<14198> A_IWL<14197> A_IWL<14196> A_IWL<14195> A_IWL<14194> A_IWL<14193> A_IWL<14192> A_IWL<14191> A_IWL<14190> A_IWL<14189> A_IWL<14188> A_IWL<14187> A_IWL<14186> A_IWL<14185> A_IWL<14184> A_IWL<14183> A_IWL<14182> A_IWL<14181> A_IWL<14180> A_IWL<14179> A_IWL<14178> A_IWL<14177> A_IWL<14176> A_IWL<14175> A_IWL<14174> A_IWL<14173> A_IWL<14172> A_IWL<14171> A_IWL<14170> A_IWL<14169> A_IWL<14168> A_IWL<14167> A_IWL<14166> A_IWL<14165> A_IWL<14164> A_IWL<14163> A_IWL<14162> A_IWL<14161> A_IWL<14160> A_IWL<14159> A_IWL<14158> A_IWL<14157> A_IWL<14156> A_IWL<14155> A_IWL<14154> A_IWL<14153> A_IWL<14152> A_IWL<14151> A_IWL<14150> A_IWL<14149> A_IWL<14148> A_IWL<14147> A_IWL<14146> A_IWL<14145> A_IWL<14144> A_IWL<14143> A_IWL<14142> A_IWL<14141> A_IWL<14140> A_IWL<14139> A_IWL<14138> A_IWL<14137> A_IWL<14136> A_IWL<14135> A_IWL<14134> A_IWL<14133> A_IWL<14132> A_IWL<14131> A_IWL<14130> A_IWL<14129> A_IWL<14128> A_IWL<14127> A_IWL<14126> A_IWL<14125> A_IWL<14124> A_IWL<14123> A_IWL<14122> A_IWL<14121> A_IWL<14120> A_IWL<14119> A_IWL<14118> A_IWL<14117> A_IWL<14116> A_IWL<14115> A_IWL<14114> A_IWL<14113> A_IWL<14112> A_IWL<14111> A_IWL<14110> A_IWL<14109> A_IWL<14108> A_IWL<14107> A_IWL<14106> A_IWL<14105> A_IWL<14104> A_IWL<14103> A_IWL<14102> A_IWL<14101> A_IWL<14100> A_IWL<14099> A_IWL<14098> A_IWL<14097> A_IWL<14096> A_IWL<14095> A_IWL<14094> A_IWL<14093> A_IWL<14092> A_IWL<14091> A_IWL<14090> A_IWL<14089> A_IWL<14088> A_IWL<14087> A_IWL<14086> A_IWL<14085> A_IWL<14084> A_IWL<14083> A_IWL<14082> A_IWL<14081> A_IWL<14080> A_IWL<14079> A_IWL<14078> A_IWL<14077> A_IWL<14076> A_IWL<14075> A_IWL<14074> A_IWL<14073> A_IWL<14072> A_IWL<14071> A_IWL<14070> A_IWL<14069> A_IWL<14068> A_IWL<14067> A_IWL<14066> A_IWL<14065> A_IWL<14064> A_IWL<14063> A_IWL<14062> A_IWL<14061> A_IWL<14060> A_IWL<14059> A_IWL<14058> A_IWL<14057> A_IWL<14056> A_IWL<14055> A_IWL<14054> A_IWL<14053> A_IWL<14052> A_IWL<14051> A_IWL<14050> A_IWL<14049> A_IWL<14048> A_IWL<14047> A_IWL<14046> A_IWL<14045> A_IWL<14044> A_IWL<14043> A_IWL<14042> A_IWL<14041> A_IWL<14040> A_IWL<14039> A_IWL<14038> A_IWL<14037> A_IWL<14036> A_IWL<14035> A_IWL<14034> A_IWL<14033> A_IWL<14032> A_IWL<14031> A_IWL<14030> A_IWL<14029> A_IWL<14028> A_IWL<14027> A_IWL<14026> A_IWL<14025> A_IWL<14024> A_IWL<14023> A_IWL<14022> A_IWL<14021> A_IWL<14020> A_IWL<14019> A_IWL<14018> A_IWL<14017> A_IWL<14016> A_IWL<14015> A_IWL<14014> A_IWL<14013> A_IWL<14012> A_IWL<14011> A_IWL<14010> A_IWL<14009> A_IWL<14008> A_IWL<14007> A_IWL<14006> A_IWL<14005> A_IWL<14004> A_IWL<14003> A_IWL<14002> A_IWL<14001> A_IWL<14000> A_IWL<13999> A_IWL<13998> A_IWL<13997> A_IWL<13996> A_IWL<13995> A_IWL<13994> A_IWL<13993> A_IWL<13992> A_IWL<13991> A_IWL<13990> A_IWL<13989> A_IWL<13988> A_IWL<13987> A_IWL<13986> A_IWL<13985> A_IWL<13984> A_IWL<13983> A_IWL<13982> A_IWL<13981> A_IWL<13980> A_IWL<13979> A_IWL<13978> A_IWL<13977> A_IWL<13976> A_IWL<13975> A_IWL<13974> A_IWL<13973> A_IWL<13972> A_IWL<13971> A_IWL<13970> A_IWL<13969> A_IWL<13968> A_IWL<13967> A_IWL<13966> A_IWL<13965> A_IWL<13964> A_IWL<13963> A_IWL<13962> A_IWL<13961> A_IWL<13960> A_IWL<13959> A_IWL<13958> A_IWL<13957> A_IWL<13956> A_IWL<13955> A_IWL<13954> A_IWL<13953> A_IWL<13952> A_IWL<13951> A_IWL<13950> A_IWL<13949> A_IWL<13948> A_IWL<13947> A_IWL<13946> A_IWL<13945> A_IWL<13944> A_IWL<13943> A_IWL<13942> A_IWL<13941> A_IWL<13940> A_IWL<13939> A_IWL<13938> A_IWL<13937> A_IWL<13936> A_IWL<13935> A_IWL<13934> A_IWL<13933> A_IWL<13932> A_IWL<13931> A_IWL<13930> A_IWL<13929> A_IWL<13928> A_IWL<13927> A_IWL<13926> A_IWL<13925> A_IWL<13924> A_IWL<13923> A_IWL<13922> A_IWL<13921> A_IWL<13920> A_IWL<13919> A_IWL<13918> A_IWL<13917> A_IWL<13916> A_IWL<13915> A_IWL<13914> A_IWL<13913> A_IWL<13912> A_IWL<13911> A_IWL<13910> A_IWL<13909> A_IWL<13908> A_IWL<13907> A_IWL<13906> A_IWL<13905> A_IWL<13904> A_IWL<13903> A_IWL<13902> A_IWL<13901> A_IWL<13900> A_IWL<13899> A_IWL<13898> A_IWL<13897> A_IWL<13896> A_IWL<13895> A_IWL<13894> A_IWL<13893> A_IWL<13892> A_IWL<13891> A_IWL<13890> A_IWL<13889> A_IWL<13888> A_IWL<13887> A_IWL<13886> A_IWL<13885> A_IWL<13884> A_IWL<13883> A_IWL<13882> A_IWL<13881> A_IWL<13880> A_IWL<13879> A_IWL<13878> A_IWL<13877> A_IWL<13876> A_IWL<13875> A_IWL<13874> A_IWL<13873> A_IWL<13872> A_IWL<13871> A_IWL<13870> A_IWL<13869> A_IWL<13868> A_IWL<13867> A_IWL<13866> A_IWL<13865> A_IWL<13864> A_IWL<13863> A_IWL<13862> A_IWL<13861> A_IWL<13860> A_IWL<13859> A_IWL<13858> A_IWL<13857> A_IWL<13856> A_IWL<13855> A_IWL<13854> A_IWL<13853> A_IWL<13852> A_IWL<13851> A_IWL<13850> A_IWL<13849> A_IWL<13848> A_IWL<13847> A_IWL<13846> A_IWL<13845> A_IWL<13844> A_IWL<13843> A_IWL<13842> A_IWL<13841> A_IWL<13840> A_IWL<13839> A_IWL<13838> A_IWL<13837> A_IWL<13836> A_IWL<13835> A_IWL<13834> A_IWL<13833> A_IWL<13832> A_IWL<13831> A_IWL<13830> A_IWL<13829> A_IWL<13828> A_IWL<13827> A_IWL<13826> A_IWL<13825> A_IWL<13824> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<26> A_BLC<53> A_BLC<52> A_BLC_TOP<53> A_BLC_TOP<52> A_BLT<53> A_BLT<52> A_BLT_TOP<53> A_BLT_TOP<52> A_IWL<13311> A_IWL<13310> A_IWL<13309> A_IWL<13308> A_IWL<13307> A_IWL<13306> A_IWL<13305> A_IWL<13304> A_IWL<13303> A_IWL<13302> A_IWL<13301> A_IWL<13300> A_IWL<13299> A_IWL<13298> A_IWL<13297> A_IWL<13296> A_IWL<13295> A_IWL<13294> A_IWL<13293> A_IWL<13292> A_IWL<13291> A_IWL<13290> A_IWL<13289> A_IWL<13288> A_IWL<13287> A_IWL<13286> A_IWL<13285> A_IWL<13284> A_IWL<13283> A_IWL<13282> A_IWL<13281> A_IWL<13280> A_IWL<13279> A_IWL<13278> A_IWL<13277> A_IWL<13276> A_IWL<13275> A_IWL<13274> A_IWL<13273> A_IWL<13272> A_IWL<13271> A_IWL<13270> A_IWL<13269> A_IWL<13268> A_IWL<13267> A_IWL<13266> A_IWL<13265> A_IWL<13264> A_IWL<13263> A_IWL<13262> A_IWL<13261> A_IWL<13260> A_IWL<13259> A_IWL<13258> A_IWL<13257> A_IWL<13256> A_IWL<13255> A_IWL<13254> A_IWL<13253> A_IWL<13252> A_IWL<13251> A_IWL<13250> A_IWL<13249> A_IWL<13248> A_IWL<13247> A_IWL<13246> A_IWL<13245> A_IWL<13244> A_IWL<13243> A_IWL<13242> A_IWL<13241> A_IWL<13240> A_IWL<13239> A_IWL<13238> A_IWL<13237> A_IWL<13236> A_IWL<13235> A_IWL<13234> A_IWL<13233> A_IWL<13232> A_IWL<13231> A_IWL<13230> A_IWL<13229> A_IWL<13228> A_IWL<13227> A_IWL<13226> A_IWL<13225> A_IWL<13224> A_IWL<13223> A_IWL<13222> A_IWL<13221> A_IWL<13220> A_IWL<13219> A_IWL<13218> A_IWL<13217> A_IWL<13216> A_IWL<13215> A_IWL<13214> A_IWL<13213> A_IWL<13212> A_IWL<13211> A_IWL<13210> A_IWL<13209> A_IWL<13208> A_IWL<13207> A_IWL<13206> A_IWL<13205> A_IWL<13204> A_IWL<13203> A_IWL<13202> A_IWL<13201> A_IWL<13200> A_IWL<13199> A_IWL<13198> A_IWL<13197> A_IWL<13196> A_IWL<13195> A_IWL<13194> A_IWL<13193> A_IWL<13192> A_IWL<13191> A_IWL<13190> A_IWL<13189> A_IWL<13188> A_IWL<13187> A_IWL<13186> A_IWL<13185> A_IWL<13184> A_IWL<13183> A_IWL<13182> A_IWL<13181> A_IWL<13180> A_IWL<13179> A_IWL<13178> A_IWL<13177> A_IWL<13176> A_IWL<13175> A_IWL<13174> A_IWL<13173> A_IWL<13172> A_IWL<13171> A_IWL<13170> A_IWL<13169> A_IWL<13168> A_IWL<13167> A_IWL<13166> A_IWL<13165> A_IWL<13164> A_IWL<13163> A_IWL<13162> A_IWL<13161> A_IWL<13160> A_IWL<13159> A_IWL<13158> A_IWL<13157> A_IWL<13156> A_IWL<13155> A_IWL<13154> A_IWL<13153> A_IWL<13152> A_IWL<13151> A_IWL<13150> A_IWL<13149> A_IWL<13148> A_IWL<13147> A_IWL<13146> A_IWL<13145> A_IWL<13144> A_IWL<13143> A_IWL<13142> A_IWL<13141> A_IWL<13140> A_IWL<13139> A_IWL<13138> A_IWL<13137> A_IWL<13136> A_IWL<13135> A_IWL<13134> A_IWL<13133> A_IWL<13132> A_IWL<13131> A_IWL<13130> A_IWL<13129> A_IWL<13128> A_IWL<13127> A_IWL<13126> A_IWL<13125> A_IWL<13124> A_IWL<13123> A_IWL<13122> A_IWL<13121> A_IWL<13120> A_IWL<13119> A_IWL<13118> A_IWL<13117> A_IWL<13116> A_IWL<13115> A_IWL<13114> A_IWL<13113> A_IWL<13112> A_IWL<13111> A_IWL<13110> A_IWL<13109> A_IWL<13108> A_IWL<13107> A_IWL<13106> A_IWL<13105> A_IWL<13104> A_IWL<13103> A_IWL<13102> A_IWL<13101> A_IWL<13100> A_IWL<13099> A_IWL<13098> A_IWL<13097> A_IWL<13096> A_IWL<13095> A_IWL<13094> A_IWL<13093> A_IWL<13092> A_IWL<13091> A_IWL<13090> A_IWL<13089> A_IWL<13088> A_IWL<13087> A_IWL<13086> A_IWL<13085> A_IWL<13084> A_IWL<13083> A_IWL<13082> A_IWL<13081> A_IWL<13080> A_IWL<13079> A_IWL<13078> A_IWL<13077> A_IWL<13076> A_IWL<13075> A_IWL<13074> A_IWL<13073> A_IWL<13072> A_IWL<13071> A_IWL<13070> A_IWL<13069> A_IWL<13068> A_IWL<13067> A_IWL<13066> A_IWL<13065> A_IWL<13064> A_IWL<13063> A_IWL<13062> A_IWL<13061> A_IWL<13060> A_IWL<13059> A_IWL<13058> A_IWL<13057> A_IWL<13056> A_IWL<13055> A_IWL<13054> A_IWL<13053> A_IWL<13052> A_IWL<13051> A_IWL<13050> A_IWL<13049> A_IWL<13048> A_IWL<13047> A_IWL<13046> A_IWL<13045> A_IWL<13044> A_IWL<13043> A_IWL<13042> A_IWL<13041> A_IWL<13040> A_IWL<13039> A_IWL<13038> A_IWL<13037> A_IWL<13036> A_IWL<13035> A_IWL<13034> A_IWL<13033> A_IWL<13032> A_IWL<13031> A_IWL<13030> A_IWL<13029> A_IWL<13028> A_IWL<13027> A_IWL<13026> A_IWL<13025> A_IWL<13024> A_IWL<13023> A_IWL<13022> A_IWL<13021> A_IWL<13020> A_IWL<13019> A_IWL<13018> A_IWL<13017> A_IWL<13016> A_IWL<13015> A_IWL<13014> A_IWL<13013> A_IWL<13012> A_IWL<13011> A_IWL<13010> A_IWL<13009> A_IWL<13008> A_IWL<13007> A_IWL<13006> A_IWL<13005> A_IWL<13004> A_IWL<13003> A_IWL<13002> A_IWL<13001> A_IWL<13000> A_IWL<12999> A_IWL<12998> A_IWL<12997> A_IWL<12996> A_IWL<12995> A_IWL<12994> A_IWL<12993> A_IWL<12992> A_IWL<12991> A_IWL<12990> A_IWL<12989> A_IWL<12988> A_IWL<12987> A_IWL<12986> A_IWL<12985> A_IWL<12984> A_IWL<12983> A_IWL<12982> A_IWL<12981> A_IWL<12980> A_IWL<12979> A_IWL<12978> A_IWL<12977> A_IWL<12976> A_IWL<12975> A_IWL<12974> A_IWL<12973> A_IWL<12972> A_IWL<12971> A_IWL<12970> A_IWL<12969> A_IWL<12968> A_IWL<12967> A_IWL<12966> A_IWL<12965> A_IWL<12964> A_IWL<12963> A_IWL<12962> A_IWL<12961> A_IWL<12960> A_IWL<12959> A_IWL<12958> A_IWL<12957> A_IWL<12956> A_IWL<12955> A_IWL<12954> A_IWL<12953> A_IWL<12952> A_IWL<12951> A_IWL<12950> A_IWL<12949> A_IWL<12948> A_IWL<12947> A_IWL<12946> A_IWL<12945> A_IWL<12944> A_IWL<12943> A_IWL<12942> A_IWL<12941> A_IWL<12940> A_IWL<12939> A_IWL<12938> A_IWL<12937> A_IWL<12936> A_IWL<12935> A_IWL<12934> A_IWL<12933> A_IWL<12932> A_IWL<12931> A_IWL<12930> A_IWL<12929> A_IWL<12928> A_IWL<12927> A_IWL<12926> A_IWL<12925> A_IWL<12924> A_IWL<12923> A_IWL<12922> A_IWL<12921> A_IWL<12920> A_IWL<12919> A_IWL<12918> A_IWL<12917> A_IWL<12916> A_IWL<12915> A_IWL<12914> A_IWL<12913> A_IWL<12912> A_IWL<12911> A_IWL<12910> A_IWL<12909> A_IWL<12908> A_IWL<12907> A_IWL<12906> A_IWL<12905> A_IWL<12904> A_IWL<12903> A_IWL<12902> A_IWL<12901> A_IWL<12900> A_IWL<12899> A_IWL<12898> A_IWL<12897> A_IWL<12896> A_IWL<12895> A_IWL<12894> A_IWL<12893> A_IWL<12892> A_IWL<12891> A_IWL<12890> A_IWL<12889> A_IWL<12888> A_IWL<12887> A_IWL<12886> A_IWL<12885> A_IWL<12884> A_IWL<12883> A_IWL<12882> A_IWL<12881> A_IWL<12880> A_IWL<12879> A_IWL<12878> A_IWL<12877> A_IWL<12876> A_IWL<12875> A_IWL<12874> A_IWL<12873> A_IWL<12872> A_IWL<12871> A_IWL<12870> A_IWL<12869> A_IWL<12868> A_IWL<12867> A_IWL<12866> A_IWL<12865> A_IWL<12864> A_IWL<12863> A_IWL<12862> A_IWL<12861> A_IWL<12860> A_IWL<12859> A_IWL<12858> A_IWL<12857> A_IWL<12856> A_IWL<12855> A_IWL<12854> A_IWL<12853> A_IWL<12852> A_IWL<12851> A_IWL<12850> A_IWL<12849> A_IWL<12848> A_IWL<12847> A_IWL<12846> A_IWL<12845> A_IWL<12844> A_IWL<12843> A_IWL<12842> A_IWL<12841> A_IWL<12840> A_IWL<12839> A_IWL<12838> A_IWL<12837> A_IWL<12836> A_IWL<12835> A_IWL<12834> A_IWL<12833> A_IWL<12832> A_IWL<12831> A_IWL<12830> A_IWL<12829> A_IWL<12828> A_IWL<12827> A_IWL<12826> A_IWL<12825> A_IWL<12824> A_IWL<12823> A_IWL<12822> A_IWL<12821> A_IWL<12820> A_IWL<12819> A_IWL<12818> A_IWL<12817> A_IWL<12816> A_IWL<12815> A_IWL<12814> A_IWL<12813> A_IWL<12812> A_IWL<12811> A_IWL<12810> A_IWL<12809> A_IWL<12808> A_IWL<12807> A_IWL<12806> A_IWL<12805> A_IWL<12804> A_IWL<12803> A_IWL<12802> A_IWL<12801> A_IWL<12800> A_IWL<13823> A_IWL<13822> A_IWL<13821> A_IWL<13820> A_IWL<13819> A_IWL<13818> A_IWL<13817> A_IWL<13816> A_IWL<13815> A_IWL<13814> A_IWL<13813> A_IWL<13812> A_IWL<13811> A_IWL<13810> A_IWL<13809> A_IWL<13808> A_IWL<13807> A_IWL<13806> A_IWL<13805> A_IWL<13804> A_IWL<13803> A_IWL<13802> A_IWL<13801> A_IWL<13800> A_IWL<13799> A_IWL<13798> A_IWL<13797> A_IWL<13796> A_IWL<13795> A_IWL<13794> A_IWL<13793> A_IWL<13792> A_IWL<13791> A_IWL<13790> A_IWL<13789> A_IWL<13788> A_IWL<13787> A_IWL<13786> A_IWL<13785> A_IWL<13784> A_IWL<13783> A_IWL<13782> A_IWL<13781> A_IWL<13780> A_IWL<13779> A_IWL<13778> A_IWL<13777> A_IWL<13776> A_IWL<13775> A_IWL<13774> A_IWL<13773> A_IWL<13772> A_IWL<13771> A_IWL<13770> A_IWL<13769> A_IWL<13768> A_IWL<13767> A_IWL<13766> A_IWL<13765> A_IWL<13764> A_IWL<13763> A_IWL<13762> A_IWL<13761> A_IWL<13760> A_IWL<13759> A_IWL<13758> A_IWL<13757> A_IWL<13756> A_IWL<13755> A_IWL<13754> A_IWL<13753> A_IWL<13752> A_IWL<13751> A_IWL<13750> A_IWL<13749> A_IWL<13748> A_IWL<13747> A_IWL<13746> A_IWL<13745> A_IWL<13744> A_IWL<13743> A_IWL<13742> A_IWL<13741> A_IWL<13740> A_IWL<13739> A_IWL<13738> A_IWL<13737> A_IWL<13736> A_IWL<13735> A_IWL<13734> A_IWL<13733> A_IWL<13732> A_IWL<13731> A_IWL<13730> A_IWL<13729> A_IWL<13728> A_IWL<13727> A_IWL<13726> A_IWL<13725> A_IWL<13724> A_IWL<13723> A_IWL<13722> A_IWL<13721> A_IWL<13720> A_IWL<13719> A_IWL<13718> A_IWL<13717> A_IWL<13716> A_IWL<13715> A_IWL<13714> A_IWL<13713> A_IWL<13712> A_IWL<13711> A_IWL<13710> A_IWL<13709> A_IWL<13708> A_IWL<13707> A_IWL<13706> A_IWL<13705> A_IWL<13704> A_IWL<13703> A_IWL<13702> A_IWL<13701> A_IWL<13700> A_IWL<13699> A_IWL<13698> A_IWL<13697> A_IWL<13696> A_IWL<13695> A_IWL<13694> A_IWL<13693> A_IWL<13692> A_IWL<13691> A_IWL<13690> A_IWL<13689> A_IWL<13688> A_IWL<13687> A_IWL<13686> A_IWL<13685> A_IWL<13684> A_IWL<13683> A_IWL<13682> A_IWL<13681> A_IWL<13680> A_IWL<13679> A_IWL<13678> A_IWL<13677> A_IWL<13676> A_IWL<13675> A_IWL<13674> A_IWL<13673> A_IWL<13672> A_IWL<13671> A_IWL<13670> A_IWL<13669> A_IWL<13668> A_IWL<13667> A_IWL<13666> A_IWL<13665> A_IWL<13664> A_IWL<13663> A_IWL<13662> A_IWL<13661> A_IWL<13660> A_IWL<13659> A_IWL<13658> A_IWL<13657> A_IWL<13656> A_IWL<13655> A_IWL<13654> A_IWL<13653> A_IWL<13652> A_IWL<13651> A_IWL<13650> A_IWL<13649> A_IWL<13648> A_IWL<13647> A_IWL<13646> A_IWL<13645> A_IWL<13644> A_IWL<13643> A_IWL<13642> A_IWL<13641> A_IWL<13640> A_IWL<13639> A_IWL<13638> A_IWL<13637> A_IWL<13636> A_IWL<13635> A_IWL<13634> A_IWL<13633> A_IWL<13632> A_IWL<13631> A_IWL<13630> A_IWL<13629> A_IWL<13628> A_IWL<13627> A_IWL<13626> A_IWL<13625> A_IWL<13624> A_IWL<13623> A_IWL<13622> A_IWL<13621> A_IWL<13620> A_IWL<13619> A_IWL<13618> A_IWL<13617> A_IWL<13616> A_IWL<13615> A_IWL<13614> A_IWL<13613> A_IWL<13612> A_IWL<13611> A_IWL<13610> A_IWL<13609> A_IWL<13608> A_IWL<13607> A_IWL<13606> A_IWL<13605> A_IWL<13604> A_IWL<13603> A_IWL<13602> A_IWL<13601> A_IWL<13600> A_IWL<13599> A_IWL<13598> A_IWL<13597> A_IWL<13596> A_IWL<13595> A_IWL<13594> A_IWL<13593> A_IWL<13592> A_IWL<13591> A_IWL<13590> A_IWL<13589> A_IWL<13588> A_IWL<13587> A_IWL<13586> A_IWL<13585> A_IWL<13584> A_IWL<13583> A_IWL<13582> A_IWL<13581> A_IWL<13580> A_IWL<13579> A_IWL<13578> A_IWL<13577> A_IWL<13576> A_IWL<13575> A_IWL<13574> A_IWL<13573> A_IWL<13572> A_IWL<13571> A_IWL<13570> A_IWL<13569> A_IWL<13568> A_IWL<13567> A_IWL<13566> A_IWL<13565> A_IWL<13564> A_IWL<13563> A_IWL<13562> A_IWL<13561> A_IWL<13560> A_IWL<13559> A_IWL<13558> A_IWL<13557> A_IWL<13556> A_IWL<13555> A_IWL<13554> A_IWL<13553> A_IWL<13552> A_IWL<13551> A_IWL<13550> A_IWL<13549> A_IWL<13548> A_IWL<13547> A_IWL<13546> A_IWL<13545> A_IWL<13544> A_IWL<13543> A_IWL<13542> A_IWL<13541> A_IWL<13540> A_IWL<13539> A_IWL<13538> A_IWL<13537> A_IWL<13536> A_IWL<13535> A_IWL<13534> A_IWL<13533> A_IWL<13532> A_IWL<13531> A_IWL<13530> A_IWL<13529> A_IWL<13528> A_IWL<13527> A_IWL<13526> A_IWL<13525> A_IWL<13524> A_IWL<13523> A_IWL<13522> A_IWL<13521> A_IWL<13520> A_IWL<13519> A_IWL<13518> A_IWL<13517> A_IWL<13516> A_IWL<13515> A_IWL<13514> A_IWL<13513> A_IWL<13512> A_IWL<13511> A_IWL<13510> A_IWL<13509> A_IWL<13508> A_IWL<13507> A_IWL<13506> A_IWL<13505> A_IWL<13504> A_IWL<13503> A_IWL<13502> A_IWL<13501> A_IWL<13500> A_IWL<13499> A_IWL<13498> A_IWL<13497> A_IWL<13496> A_IWL<13495> A_IWL<13494> A_IWL<13493> A_IWL<13492> A_IWL<13491> A_IWL<13490> A_IWL<13489> A_IWL<13488> A_IWL<13487> A_IWL<13486> A_IWL<13485> A_IWL<13484> A_IWL<13483> A_IWL<13482> A_IWL<13481> A_IWL<13480> A_IWL<13479> A_IWL<13478> A_IWL<13477> A_IWL<13476> A_IWL<13475> A_IWL<13474> A_IWL<13473> A_IWL<13472> A_IWL<13471> A_IWL<13470> A_IWL<13469> A_IWL<13468> A_IWL<13467> A_IWL<13466> A_IWL<13465> A_IWL<13464> A_IWL<13463> A_IWL<13462> A_IWL<13461> A_IWL<13460> A_IWL<13459> A_IWL<13458> A_IWL<13457> A_IWL<13456> A_IWL<13455> A_IWL<13454> A_IWL<13453> A_IWL<13452> A_IWL<13451> A_IWL<13450> A_IWL<13449> A_IWL<13448> A_IWL<13447> A_IWL<13446> A_IWL<13445> A_IWL<13444> A_IWL<13443> A_IWL<13442> A_IWL<13441> A_IWL<13440> A_IWL<13439> A_IWL<13438> A_IWL<13437> A_IWL<13436> A_IWL<13435> A_IWL<13434> A_IWL<13433> A_IWL<13432> A_IWL<13431> A_IWL<13430> A_IWL<13429> A_IWL<13428> A_IWL<13427> A_IWL<13426> A_IWL<13425> A_IWL<13424> A_IWL<13423> A_IWL<13422> A_IWL<13421> A_IWL<13420> A_IWL<13419> A_IWL<13418> A_IWL<13417> A_IWL<13416> A_IWL<13415> A_IWL<13414> A_IWL<13413> A_IWL<13412> A_IWL<13411> A_IWL<13410> A_IWL<13409> A_IWL<13408> A_IWL<13407> A_IWL<13406> A_IWL<13405> A_IWL<13404> A_IWL<13403> A_IWL<13402> A_IWL<13401> A_IWL<13400> A_IWL<13399> A_IWL<13398> A_IWL<13397> A_IWL<13396> A_IWL<13395> A_IWL<13394> A_IWL<13393> A_IWL<13392> A_IWL<13391> A_IWL<13390> A_IWL<13389> A_IWL<13388> A_IWL<13387> A_IWL<13386> A_IWL<13385> A_IWL<13384> A_IWL<13383> A_IWL<13382> A_IWL<13381> A_IWL<13380> A_IWL<13379> A_IWL<13378> A_IWL<13377> A_IWL<13376> A_IWL<13375> A_IWL<13374> A_IWL<13373> A_IWL<13372> A_IWL<13371> A_IWL<13370> A_IWL<13369> A_IWL<13368> A_IWL<13367> A_IWL<13366> A_IWL<13365> A_IWL<13364> A_IWL<13363> A_IWL<13362> A_IWL<13361> A_IWL<13360> A_IWL<13359> A_IWL<13358> A_IWL<13357> A_IWL<13356> A_IWL<13355> A_IWL<13354> A_IWL<13353> A_IWL<13352> A_IWL<13351> A_IWL<13350> A_IWL<13349> A_IWL<13348> A_IWL<13347> A_IWL<13346> A_IWL<13345> A_IWL<13344> A_IWL<13343> A_IWL<13342> A_IWL<13341> A_IWL<13340> A_IWL<13339> A_IWL<13338> A_IWL<13337> A_IWL<13336> A_IWL<13335> A_IWL<13334> A_IWL<13333> A_IWL<13332> A_IWL<13331> A_IWL<13330> A_IWL<13329> A_IWL<13328> A_IWL<13327> A_IWL<13326> A_IWL<13325> A_IWL<13324> A_IWL<13323> A_IWL<13322> A_IWL<13321> A_IWL<13320> A_IWL<13319> A_IWL<13318> A_IWL<13317> A_IWL<13316> A_IWL<13315> A_IWL<13314> A_IWL<13313> A_IWL<13312> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<25> A_BLC<51> A_BLC<50> A_BLC_TOP<51> A_BLC_TOP<50> A_BLT<51> A_BLT<50> A_BLT_TOP<51> A_BLT_TOP<50> A_IWL<12799> A_IWL<12798> A_IWL<12797> A_IWL<12796> A_IWL<12795> A_IWL<12794> A_IWL<12793> A_IWL<12792> A_IWL<12791> A_IWL<12790> A_IWL<12789> A_IWL<12788> A_IWL<12787> A_IWL<12786> A_IWL<12785> A_IWL<12784> A_IWL<12783> A_IWL<12782> A_IWL<12781> A_IWL<12780> A_IWL<12779> A_IWL<12778> A_IWL<12777> A_IWL<12776> A_IWL<12775> A_IWL<12774> A_IWL<12773> A_IWL<12772> A_IWL<12771> A_IWL<12770> A_IWL<12769> A_IWL<12768> A_IWL<12767> A_IWL<12766> A_IWL<12765> A_IWL<12764> A_IWL<12763> A_IWL<12762> A_IWL<12761> A_IWL<12760> A_IWL<12759> A_IWL<12758> A_IWL<12757> A_IWL<12756> A_IWL<12755> A_IWL<12754> A_IWL<12753> A_IWL<12752> A_IWL<12751> A_IWL<12750> A_IWL<12749> A_IWL<12748> A_IWL<12747> A_IWL<12746> A_IWL<12745> A_IWL<12744> A_IWL<12743> A_IWL<12742> A_IWL<12741> A_IWL<12740> A_IWL<12739> A_IWL<12738> A_IWL<12737> A_IWL<12736> A_IWL<12735> A_IWL<12734> A_IWL<12733> A_IWL<12732> A_IWL<12731> A_IWL<12730> A_IWL<12729> A_IWL<12728> A_IWL<12727> A_IWL<12726> A_IWL<12725> A_IWL<12724> A_IWL<12723> A_IWL<12722> A_IWL<12721> A_IWL<12720> A_IWL<12719> A_IWL<12718> A_IWL<12717> A_IWL<12716> A_IWL<12715> A_IWL<12714> A_IWL<12713> A_IWL<12712> A_IWL<12711> A_IWL<12710> A_IWL<12709> A_IWL<12708> A_IWL<12707> A_IWL<12706> A_IWL<12705> A_IWL<12704> A_IWL<12703> A_IWL<12702> A_IWL<12701> A_IWL<12700> A_IWL<12699> A_IWL<12698> A_IWL<12697> A_IWL<12696> A_IWL<12695> A_IWL<12694> A_IWL<12693> A_IWL<12692> A_IWL<12691> A_IWL<12690> A_IWL<12689> A_IWL<12688> A_IWL<12687> A_IWL<12686> A_IWL<12685> A_IWL<12684> A_IWL<12683> A_IWL<12682> A_IWL<12681> A_IWL<12680> A_IWL<12679> A_IWL<12678> A_IWL<12677> A_IWL<12676> A_IWL<12675> A_IWL<12674> A_IWL<12673> A_IWL<12672> A_IWL<12671> A_IWL<12670> A_IWL<12669> A_IWL<12668> A_IWL<12667> A_IWL<12666> A_IWL<12665> A_IWL<12664> A_IWL<12663> A_IWL<12662> A_IWL<12661> A_IWL<12660> A_IWL<12659> A_IWL<12658> A_IWL<12657> A_IWL<12656> A_IWL<12655> A_IWL<12654> A_IWL<12653> A_IWL<12652> A_IWL<12651> A_IWL<12650> A_IWL<12649> A_IWL<12648> A_IWL<12647> A_IWL<12646> A_IWL<12645> A_IWL<12644> A_IWL<12643> A_IWL<12642> A_IWL<12641> A_IWL<12640> A_IWL<12639> A_IWL<12638> A_IWL<12637> A_IWL<12636> A_IWL<12635> A_IWL<12634> A_IWL<12633> A_IWL<12632> A_IWL<12631> A_IWL<12630> A_IWL<12629> A_IWL<12628> A_IWL<12627> A_IWL<12626> A_IWL<12625> A_IWL<12624> A_IWL<12623> A_IWL<12622> A_IWL<12621> A_IWL<12620> A_IWL<12619> A_IWL<12618> A_IWL<12617> A_IWL<12616> A_IWL<12615> A_IWL<12614> A_IWL<12613> A_IWL<12612> A_IWL<12611> A_IWL<12610> A_IWL<12609> A_IWL<12608> A_IWL<12607> A_IWL<12606> A_IWL<12605> A_IWL<12604> A_IWL<12603> A_IWL<12602> A_IWL<12601> A_IWL<12600> A_IWL<12599> A_IWL<12598> A_IWL<12597> A_IWL<12596> A_IWL<12595> A_IWL<12594> A_IWL<12593> A_IWL<12592> A_IWL<12591> A_IWL<12590> A_IWL<12589> A_IWL<12588> A_IWL<12587> A_IWL<12586> A_IWL<12585> A_IWL<12584> A_IWL<12583> A_IWL<12582> A_IWL<12581> A_IWL<12580> A_IWL<12579> A_IWL<12578> A_IWL<12577> A_IWL<12576> A_IWL<12575> A_IWL<12574> A_IWL<12573> A_IWL<12572> A_IWL<12571> A_IWL<12570> A_IWL<12569> A_IWL<12568> A_IWL<12567> A_IWL<12566> A_IWL<12565> A_IWL<12564> A_IWL<12563> A_IWL<12562> A_IWL<12561> A_IWL<12560> A_IWL<12559> A_IWL<12558> A_IWL<12557> A_IWL<12556> A_IWL<12555> A_IWL<12554> A_IWL<12553> A_IWL<12552> A_IWL<12551> A_IWL<12550> A_IWL<12549> A_IWL<12548> A_IWL<12547> A_IWL<12546> A_IWL<12545> A_IWL<12544> A_IWL<12543> A_IWL<12542> A_IWL<12541> A_IWL<12540> A_IWL<12539> A_IWL<12538> A_IWL<12537> A_IWL<12536> A_IWL<12535> A_IWL<12534> A_IWL<12533> A_IWL<12532> A_IWL<12531> A_IWL<12530> A_IWL<12529> A_IWL<12528> A_IWL<12527> A_IWL<12526> A_IWL<12525> A_IWL<12524> A_IWL<12523> A_IWL<12522> A_IWL<12521> A_IWL<12520> A_IWL<12519> A_IWL<12518> A_IWL<12517> A_IWL<12516> A_IWL<12515> A_IWL<12514> A_IWL<12513> A_IWL<12512> A_IWL<12511> A_IWL<12510> A_IWL<12509> A_IWL<12508> A_IWL<12507> A_IWL<12506> A_IWL<12505> A_IWL<12504> A_IWL<12503> A_IWL<12502> A_IWL<12501> A_IWL<12500> A_IWL<12499> A_IWL<12498> A_IWL<12497> A_IWL<12496> A_IWL<12495> A_IWL<12494> A_IWL<12493> A_IWL<12492> A_IWL<12491> A_IWL<12490> A_IWL<12489> A_IWL<12488> A_IWL<12487> A_IWL<12486> A_IWL<12485> A_IWL<12484> A_IWL<12483> A_IWL<12482> A_IWL<12481> A_IWL<12480> A_IWL<12479> A_IWL<12478> A_IWL<12477> A_IWL<12476> A_IWL<12475> A_IWL<12474> A_IWL<12473> A_IWL<12472> A_IWL<12471> A_IWL<12470> A_IWL<12469> A_IWL<12468> A_IWL<12467> A_IWL<12466> A_IWL<12465> A_IWL<12464> A_IWL<12463> A_IWL<12462> A_IWL<12461> A_IWL<12460> A_IWL<12459> A_IWL<12458> A_IWL<12457> A_IWL<12456> A_IWL<12455> A_IWL<12454> A_IWL<12453> A_IWL<12452> A_IWL<12451> A_IWL<12450> A_IWL<12449> A_IWL<12448> A_IWL<12447> A_IWL<12446> A_IWL<12445> A_IWL<12444> A_IWL<12443> A_IWL<12442> A_IWL<12441> A_IWL<12440> A_IWL<12439> A_IWL<12438> A_IWL<12437> A_IWL<12436> A_IWL<12435> A_IWL<12434> A_IWL<12433> A_IWL<12432> A_IWL<12431> A_IWL<12430> A_IWL<12429> A_IWL<12428> A_IWL<12427> A_IWL<12426> A_IWL<12425> A_IWL<12424> A_IWL<12423> A_IWL<12422> A_IWL<12421> A_IWL<12420> A_IWL<12419> A_IWL<12418> A_IWL<12417> A_IWL<12416> A_IWL<12415> A_IWL<12414> A_IWL<12413> A_IWL<12412> A_IWL<12411> A_IWL<12410> A_IWL<12409> A_IWL<12408> A_IWL<12407> A_IWL<12406> A_IWL<12405> A_IWL<12404> A_IWL<12403> A_IWL<12402> A_IWL<12401> A_IWL<12400> A_IWL<12399> A_IWL<12398> A_IWL<12397> A_IWL<12396> A_IWL<12395> A_IWL<12394> A_IWL<12393> A_IWL<12392> A_IWL<12391> A_IWL<12390> A_IWL<12389> A_IWL<12388> A_IWL<12387> A_IWL<12386> A_IWL<12385> A_IWL<12384> A_IWL<12383> A_IWL<12382> A_IWL<12381> A_IWL<12380> A_IWL<12379> A_IWL<12378> A_IWL<12377> A_IWL<12376> A_IWL<12375> A_IWL<12374> A_IWL<12373> A_IWL<12372> A_IWL<12371> A_IWL<12370> A_IWL<12369> A_IWL<12368> A_IWL<12367> A_IWL<12366> A_IWL<12365> A_IWL<12364> A_IWL<12363> A_IWL<12362> A_IWL<12361> A_IWL<12360> A_IWL<12359> A_IWL<12358> A_IWL<12357> A_IWL<12356> A_IWL<12355> A_IWL<12354> A_IWL<12353> A_IWL<12352> A_IWL<12351> A_IWL<12350> A_IWL<12349> A_IWL<12348> A_IWL<12347> A_IWL<12346> A_IWL<12345> A_IWL<12344> A_IWL<12343> A_IWL<12342> A_IWL<12341> A_IWL<12340> A_IWL<12339> A_IWL<12338> A_IWL<12337> A_IWL<12336> A_IWL<12335> A_IWL<12334> A_IWL<12333> A_IWL<12332> A_IWL<12331> A_IWL<12330> A_IWL<12329> A_IWL<12328> A_IWL<12327> A_IWL<12326> A_IWL<12325> A_IWL<12324> A_IWL<12323> A_IWL<12322> A_IWL<12321> A_IWL<12320> A_IWL<12319> A_IWL<12318> A_IWL<12317> A_IWL<12316> A_IWL<12315> A_IWL<12314> A_IWL<12313> A_IWL<12312> A_IWL<12311> A_IWL<12310> A_IWL<12309> A_IWL<12308> A_IWL<12307> A_IWL<12306> A_IWL<12305> A_IWL<12304> A_IWL<12303> A_IWL<12302> A_IWL<12301> A_IWL<12300> A_IWL<12299> A_IWL<12298> A_IWL<12297> A_IWL<12296> A_IWL<12295> A_IWL<12294> A_IWL<12293> A_IWL<12292> A_IWL<12291> A_IWL<12290> A_IWL<12289> A_IWL<12288> A_IWL<13311> A_IWL<13310> A_IWL<13309> A_IWL<13308> A_IWL<13307> A_IWL<13306> A_IWL<13305> A_IWL<13304> A_IWL<13303> A_IWL<13302> A_IWL<13301> A_IWL<13300> A_IWL<13299> A_IWL<13298> A_IWL<13297> A_IWL<13296> A_IWL<13295> A_IWL<13294> A_IWL<13293> A_IWL<13292> A_IWL<13291> A_IWL<13290> A_IWL<13289> A_IWL<13288> A_IWL<13287> A_IWL<13286> A_IWL<13285> A_IWL<13284> A_IWL<13283> A_IWL<13282> A_IWL<13281> A_IWL<13280> A_IWL<13279> A_IWL<13278> A_IWL<13277> A_IWL<13276> A_IWL<13275> A_IWL<13274> A_IWL<13273> A_IWL<13272> A_IWL<13271> A_IWL<13270> A_IWL<13269> A_IWL<13268> A_IWL<13267> A_IWL<13266> A_IWL<13265> A_IWL<13264> A_IWL<13263> A_IWL<13262> A_IWL<13261> A_IWL<13260> A_IWL<13259> A_IWL<13258> A_IWL<13257> A_IWL<13256> A_IWL<13255> A_IWL<13254> A_IWL<13253> A_IWL<13252> A_IWL<13251> A_IWL<13250> A_IWL<13249> A_IWL<13248> A_IWL<13247> A_IWL<13246> A_IWL<13245> A_IWL<13244> A_IWL<13243> A_IWL<13242> A_IWL<13241> A_IWL<13240> A_IWL<13239> A_IWL<13238> A_IWL<13237> A_IWL<13236> A_IWL<13235> A_IWL<13234> A_IWL<13233> A_IWL<13232> A_IWL<13231> A_IWL<13230> A_IWL<13229> A_IWL<13228> A_IWL<13227> A_IWL<13226> A_IWL<13225> A_IWL<13224> A_IWL<13223> A_IWL<13222> A_IWL<13221> A_IWL<13220> A_IWL<13219> A_IWL<13218> A_IWL<13217> A_IWL<13216> A_IWL<13215> A_IWL<13214> A_IWL<13213> A_IWL<13212> A_IWL<13211> A_IWL<13210> A_IWL<13209> A_IWL<13208> A_IWL<13207> A_IWL<13206> A_IWL<13205> A_IWL<13204> A_IWL<13203> A_IWL<13202> A_IWL<13201> A_IWL<13200> A_IWL<13199> A_IWL<13198> A_IWL<13197> A_IWL<13196> A_IWL<13195> A_IWL<13194> A_IWL<13193> A_IWL<13192> A_IWL<13191> A_IWL<13190> A_IWL<13189> A_IWL<13188> A_IWL<13187> A_IWL<13186> A_IWL<13185> A_IWL<13184> A_IWL<13183> A_IWL<13182> A_IWL<13181> A_IWL<13180> A_IWL<13179> A_IWL<13178> A_IWL<13177> A_IWL<13176> A_IWL<13175> A_IWL<13174> A_IWL<13173> A_IWL<13172> A_IWL<13171> A_IWL<13170> A_IWL<13169> A_IWL<13168> A_IWL<13167> A_IWL<13166> A_IWL<13165> A_IWL<13164> A_IWL<13163> A_IWL<13162> A_IWL<13161> A_IWL<13160> A_IWL<13159> A_IWL<13158> A_IWL<13157> A_IWL<13156> A_IWL<13155> A_IWL<13154> A_IWL<13153> A_IWL<13152> A_IWL<13151> A_IWL<13150> A_IWL<13149> A_IWL<13148> A_IWL<13147> A_IWL<13146> A_IWL<13145> A_IWL<13144> A_IWL<13143> A_IWL<13142> A_IWL<13141> A_IWL<13140> A_IWL<13139> A_IWL<13138> A_IWL<13137> A_IWL<13136> A_IWL<13135> A_IWL<13134> A_IWL<13133> A_IWL<13132> A_IWL<13131> A_IWL<13130> A_IWL<13129> A_IWL<13128> A_IWL<13127> A_IWL<13126> A_IWL<13125> A_IWL<13124> A_IWL<13123> A_IWL<13122> A_IWL<13121> A_IWL<13120> A_IWL<13119> A_IWL<13118> A_IWL<13117> A_IWL<13116> A_IWL<13115> A_IWL<13114> A_IWL<13113> A_IWL<13112> A_IWL<13111> A_IWL<13110> A_IWL<13109> A_IWL<13108> A_IWL<13107> A_IWL<13106> A_IWL<13105> A_IWL<13104> A_IWL<13103> A_IWL<13102> A_IWL<13101> A_IWL<13100> A_IWL<13099> A_IWL<13098> A_IWL<13097> A_IWL<13096> A_IWL<13095> A_IWL<13094> A_IWL<13093> A_IWL<13092> A_IWL<13091> A_IWL<13090> A_IWL<13089> A_IWL<13088> A_IWL<13087> A_IWL<13086> A_IWL<13085> A_IWL<13084> A_IWL<13083> A_IWL<13082> A_IWL<13081> A_IWL<13080> A_IWL<13079> A_IWL<13078> A_IWL<13077> A_IWL<13076> A_IWL<13075> A_IWL<13074> A_IWL<13073> A_IWL<13072> A_IWL<13071> A_IWL<13070> A_IWL<13069> A_IWL<13068> A_IWL<13067> A_IWL<13066> A_IWL<13065> A_IWL<13064> A_IWL<13063> A_IWL<13062> A_IWL<13061> A_IWL<13060> A_IWL<13059> A_IWL<13058> A_IWL<13057> A_IWL<13056> A_IWL<13055> A_IWL<13054> A_IWL<13053> A_IWL<13052> A_IWL<13051> A_IWL<13050> A_IWL<13049> A_IWL<13048> A_IWL<13047> A_IWL<13046> A_IWL<13045> A_IWL<13044> A_IWL<13043> A_IWL<13042> A_IWL<13041> A_IWL<13040> A_IWL<13039> A_IWL<13038> A_IWL<13037> A_IWL<13036> A_IWL<13035> A_IWL<13034> A_IWL<13033> A_IWL<13032> A_IWL<13031> A_IWL<13030> A_IWL<13029> A_IWL<13028> A_IWL<13027> A_IWL<13026> A_IWL<13025> A_IWL<13024> A_IWL<13023> A_IWL<13022> A_IWL<13021> A_IWL<13020> A_IWL<13019> A_IWL<13018> A_IWL<13017> A_IWL<13016> A_IWL<13015> A_IWL<13014> A_IWL<13013> A_IWL<13012> A_IWL<13011> A_IWL<13010> A_IWL<13009> A_IWL<13008> A_IWL<13007> A_IWL<13006> A_IWL<13005> A_IWL<13004> A_IWL<13003> A_IWL<13002> A_IWL<13001> A_IWL<13000> A_IWL<12999> A_IWL<12998> A_IWL<12997> A_IWL<12996> A_IWL<12995> A_IWL<12994> A_IWL<12993> A_IWL<12992> A_IWL<12991> A_IWL<12990> A_IWL<12989> A_IWL<12988> A_IWL<12987> A_IWL<12986> A_IWL<12985> A_IWL<12984> A_IWL<12983> A_IWL<12982> A_IWL<12981> A_IWL<12980> A_IWL<12979> A_IWL<12978> A_IWL<12977> A_IWL<12976> A_IWL<12975> A_IWL<12974> A_IWL<12973> A_IWL<12972> A_IWL<12971> A_IWL<12970> A_IWL<12969> A_IWL<12968> A_IWL<12967> A_IWL<12966> A_IWL<12965> A_IWL<12964> A_IWL<12963> A_IWL<12962> A_IWL<12961> A_IWL<12960> A_IWL<12959> A_IWL<12958> A_IWL<12957> A_IWL<12956> A_IWL<12955> A_IWL<12954> A_IWL<12953> A_IWL<12952> A_IWL<12951> A_IWL<12950> A_IWL<12949> A_IWL<12948> A_IWL<12947> A_IWL<12946> A_IWL<12945> A_IWL<12944> A_IWL<12943> A_IWL<12942> A_IWL<12941> A_IWL<12940> A_IWL<12939> A_IWL<12938> A_IWL<12937> A_IWL<12936> A_IWL<12935> A_IWL<12934> A_IWL<12933> A_IWL<12932> A_IWL<12931> A_IWL<12930> A_IWL<12929> A_IWL<12928> A_IWL<12927> A_IWL<12926> A_IWL<12925> A_IWL<12924> A_IWL<12923> A_IWL<12922> A_IWL<12921> A_IWL<12920> A_IWL<12919> A_IWL<12918> A_IWL<12917> A_IWL<12916> A_IWL<12915> A_IWL<12914> A_IWL<12913> A_IWL<12912> A_IWL<12911> A_IWL<12910> A_IWL<12909> A_IWL<12908> A_IWL<12907> A_IWL<12906> A_IWL<12905> A_IWL<12904> A_IWL<12903> A_IWL<12902> A_IWL<12901> A_IWL<12900> A_IWL<12899> A_IWL<12898> A_IWL<12897> A_IWL<12896> A_IWL<12895> A_IWL<12894> A_IWL<12893> A_IWL<12892> A_IWL<12891> A_IWL<12890> A_IWL<12889> A_IWL<12888> A_IWL<12887> A_IWL<12886> A_IWL<12885> A_IWL<12884> A_IWL<12883> A_IWL<12882> A_IWL<12881> A_IWL<12880> A_IWL<12879> A_IWL<12878> A_IWL<12877> A_IWL<12876> A_IWL<12875> A_IWL<12874> A_IWL<12873> A_IWL<12872> A_IWL<12871> A_IWL<12870> A_IWL<12869> A_IWL<12868> A_IWL<12867> A_IWL<12866> A_IWL<12865> A_IWL<12864> A_IWL<12863> A_IWL<12862> A_IWL<12861> A_IWL<12860> A_IWL<12859> A_IWL<12858> A_IWL<12857> A_IWL<12856> A_IWL<12855> A_IWL<12854> A_IWL<12853> A_IWL<12852> A_IWL<12851> A_IWL<12850> A_IWL<12849> A_IWL<12848> A_IWL<12847> A_IWL<12846> A_IWL<12845> A_IWL<12844> A_IWL<12843> A_IWL<12842> A_IWL<12841> A_IWL<12840> A_IWL<12839> A_IWL<12838> A_IWL<12837> A_IWL<12836> A_IWL<12835> A_IWL<12834> A_IWL<12833> A_IWL<12832> A_IWL<12831> A_IWL<12830> A_IWL<12829> A_IWL<12828> A_IWL<12827> A_IWL<12826> A_IWL<12825> A_IWL<12824> A_IWL<12823> A_IWL<12822> A_IWL<12821> A_IWL<12820> A_IWL<12819> A_IWL<12818> A_IWL<12817> A_IWL<12816> A_IWL<12815> A_IWL<12814> A_IWL<12813> A_IWL<12812> A_IWL<12811> A_IWL<12810> A_IWL<12809> A_IWL<12808> A_IWL<12807> A_IWL<12806> A_IWL<12805> A_IWL<12804> A_IWL<12803> A_IWL<12802> A_IWL<12801> A_IWL<12800> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<24> A_BLC<49> A_BLC<48> A_BLC_TOP<49> A_BLC_TOP<48> A_BLT<49> A_BLT<48> A_BLT_TOP<49> A_BLT_TOP<48> A_IWL<12287> A_IWL<12286> A_IWL<12285> A_IWL<12284> A_IWL<12283> A_IWL<12282> A_IWL<12281> A_IWL<12280> A_IWL<12279> A_IWL<12278> A_IWL<12277> A_IWL<12276> A_IWL<12275> A_IWL<12274> A_IWL<12273> A_IWL<12272> A_IWL<12271> A_IWL<12270> A_IWL<12269> A_IWL<12268> A_IWL<12267> A_IWL<12266> A_IWL<12265> A_IWL<12264> A_IWL<12263> A_IWL<12262> A_IWL<12261> A_IWL<12260> A_IWL<12259> A_IWL<12258> A_IWL<12257> A_IWL<12256> A_IWL<12255> A_IWL<12254> A_IWL<12253> A_IWL<12252> A_IWL<12251> A_IWL<12250> A_IWL<12249> A_IWL<12248> A_IWL<12247> A_IWL<12246> A_IWL<12245> A_IWL<12244> A_IWL<12243> A_IWL<12242> A_IWL<12241> A_IWL<12240> A_IWL<12239> A_IWL<12238> A_IWL<12237> A_IWL<12236> A_IWL<12235> A_IWL<12234> A_IWL<12233> A_IWL<12232> A_IWL<12231> A_IWL<12230> A_IWL<12229> A_IWL<12228> A_IWL<12227> A_IWL<12226> A_IWL<12225> A_IWL<12224> A_IWL<12223> A_IWL<12222> A_IWL<12221> A_IWL<12220> A_IWL<12219> A_IWL<12218> A_IWL<12217> A_IWL<12216> A_IWL<12215> A_IWL<12214> A_IWL<12213> A_IWL<12212> A_IWL<12211> A_IWL<12210> A_IWL<12209> A_IWL<12208> A_IWL<12207> A_IWL<12206> A_IWL<12205> A_IWL<12204> A_IWL<12203> A_IWL<12202> A_IWL<12201> A_IWL<12200> A_IWL<12199> A_IWL<12198> A_IWL<12197> A_IWL<12196> A_IWL<12195> A_IWL<12194> A_IWL<12193> A_IWL<12192> A_IWL<12191> A_IWL<12190> A_IWL<12189> A_IWL<12188> A_IWL<12187> A_IWL<12186> A_IWL<12185> A_IWL<12184> A_IWL<12183> A_IWL<12182> A_IWL<12181> A_IWL<12180> A_IWL<12179> A_IWL<12178> A_IWL<12177> A_IWL<12176> A_IWL<12175> A_IWL<12174> A_IWL<12173> A_IWL<12172> A_IWL<12171> A_IWL<12170> A_IWL<12169> A_IWL<12168> A_IWL<12167> A_IWL<12166> A_IWL<12165> A_IWL<12164> A_IWL<12163> A_IWL<12162> A_IWL<12161> A_IWL<12160> A_IWL<12159> A_IWL<12158> A_IWL<12157> A_IWL<12156> A_IWL<12155> A_IWL<12154> A_IWL<12153> A_IWL<12152> A_IWL<12151> A_IWL<12150> A_IWL<12149> A_IWL<12148> A_IWL<12147> A_IWL<12146> A_IWL<12145> A_IWL<12144> A_IWL<12143> A_IWL<12142> A_IWL<12141> A_IWL<12140> A_IWL<12139> A_IWL<12138> A_IWL<12137> A_IWL<12136> A_IWL<12135> A_IWL<12134> A_IWL<12133> A_IWL<12132> A_IWL<12131> A_IWL<12130> A_IWL<12129> A_IWL<12128> A_IWL<12127> A_IWL<12126> A_IWL<12125> A_IWL<12124> A_IWL<12123> A_IWL<12122> A_IWL<12121> A_IWL<12120> A_IWL<12119> A_IWL<12118> A_IWL<12117> A_IWL<12116> A_IWL<12115> A_IWL<12114> A_IWL<12113> A_IWL<12112> A_IWL<12111> A_IWL<12110> A_IWL<12109> A_IWL<12108> A_IWL<12107> A_IWL<12106> A_IWL<12105> A_IWL<12104> A_IWL<12103> A_IWL<12102> A_IWL<12101> A_IWL<12100> A_IWL<12099> A_IWL<12098> A_IWL<12097> A_IWL<12096> A_IWL<12095> A_IWL<12094> A_IWL<12093> A_IWL<12092> A_IWL<12091> A_IWL<12090> A_IWL<12089> A_IWL<12088> A_IWL<12087> A_IWL<12086> A_IWL<12085> A_IWL<12084> A_IWL<12083> A_IWL<12082> A_IWL<12081> A_IWL<12080> A_IWL<12079> A_IWL<12078> A_IWL<12077> A_IWL<12076> A_IWL<12075> A_IWL<12074> A_IWL<12073> A_IWL<12072> A_IWL<12071> A_IWL<12070> A_IWL<12069> A_IWL<12068> A_IWL<12067> A_IWL<12066> A_IWL<12065> A_IWL<12064> A_IWL<12063> A_IWL<12062> A_IWL<12061> A_IWL<12060> A_IWL<12059> A_IWL<12058> A_IWL<12057> A_IWL<12056> A_IWL<12055> A_IWL<12054> A_IWL<12053> A_IWL<12052> A_IWL<12051> A_IWL<12050> A_IWL<12049> A_IWL<12048> A_IWL<12047> A_IWL<12046> A_IWL<12045> A_IWL<12044> A_IWL<12043> A_IWL<12042> A_IWL<12041> A_IWL<12040> A_IWL<12039> A_IWL<12038> A_IWL<12037> A_IWL<12036> A_IWL<12035> A_IWL<12034> A_IWL<12033> A_IWL<12032> A_IWL<12031> A_IWL<12030> A_IWL<12029> A_IWL<12028> A_IWL<12027> A_IWL<12026> A_IWL<12025> A_IWL<12024> A_IWL<12023> A_IWL<12022> A_IWL<12021> A_IWL<12020> A_IWL<12019> A_IWL<12018> A_IWL<12017> A_IWL<12016> A_IWL<12015> A_IWL<12014> A_IWL<12013> A_IWL<12012> A_IWL<12011> A_IWL<12010> A_IWL<12009> A_IWL<12008> A_IWL<12007> A_IWL<12006> A_IWL<12005> A_IWL<12004> A_IWL<12003> A_IWL<12002> A_IWL<12001> A_IWL<12000> A_IWL<11999> A_IWL<11998> A_IWL<11997> A_IWL<11996> A_IWL<11995> A_IWL<11994> A_IWL<11993> A_IWL<11992> A_IWL<11991> A_IWL<11990> A_IWL<11989> A_IWL<11988> A_IWL<11987> A_IWL<11986> A_IWL<11985> A_IWL<11984> A_IWL<11983> A_IWL<11982> A_IWL<11981> A_IWL<11980> A_IWL<11979> A_IWL<11978> A_IWL<11977> A_IWL<11976> A_IWL<11975> A_IWL<11974> A_IWL<11973> A_IWL<11972> A_IWL<11971> A_IWL<11970> A_IWL<11969> A_IWL<11968> A_IWL<11967> A_IWL<11966> A_IWL<11965> A_IWL<11964> A_IWL<11963> A_IWL<11962> A_IWL<11961> A_IWL<11960> A_IWL<11959> A_IWL<11958> A_IWL<11957> A_IWL<11956> A_IWL<11955> A_IWL<11954> A_IWL<11953> A_IWL<11952> A_IWL<11951> A_IWL<11950> A_IWL<11949> A_IWL<11948> A_IWL<11947> A_IWL<11946> A_IWL<11945> A_IWL<11944> A_IWL<11943> A_IWL<11942> A_IWL<11941> A_IWL<11940> A_IWL<11939> A_IWL<11938> A_IWL<11937> A_IWL<11936> A_IWL<11935> A_IWL<11934> A_IWL<11933> A_IWL<11932> A_IWL<11931> A_IWL<11930> A_IWL<11929> A_IWL<11928> A_IWL<11927> A_IWL<11926> A_IWL<11925> A_IWL<11924> A_IWL<11923> A_IWL<11922> A_IWL<11921> A_IWL<11920> A_IWL<11919> A_IWL<11918> A_IWL<11917> A_IWL<11916> A_IWL<11915> A_IWL<11914> A_IWL<11913> A_IWL<11912> A_IWL<11911> A_IWL<11910> A_IWL<11909> A_IWL<11908> A_IWL<11907> A_IWL<11906> A_IWL<11905> A_IWL<11904> A_IWL<11903> A_IWL<11902> A_IWL<11901> A_IWL<11900> A_IWL<11899> A_IWL<11898> A_IWL<11897> A_IWL<11896> A_IWL<11895> A_IWL<11894> A_IWL<11893> A_IWL<11892> A_IWL<11891> A_IWL<11890> A_IWL<11889> A_IWL<11888> A_IWL<11887> A_IWL<11886> A_IWL<11885> A_IWL<11884> A_IWL<11883> A_IWL<11882> A_IWL<11881> A_IWL<11880> A_IWL<11879> A_IWL<11878> A_IWL<11877> A_IWL<11876> A_IWL<11875> A_IWL<11874> A_IWL<11873> A_IWL<11872> A_IWL<11871> A_IWL<11870> A_IWL<11869> A_IWL<11868> A_IWL<11867> A_IWL<11866> A_IWL<11865> A_IWL<11864> A_IWL<11863> A_IWL<11862> A_IWL<11861> A_IWL<11860> A_IWL<11859> A_IWL<11858> A_IWL<11857> A_IWL<11856> A_IWL<11855> A_IWL<11854> A_IWL<11853> A_IWL<11852> A_IWL<11851> A_IWL<11850> A_IWL<11849> A_IWL<11848> A_IWL<11847> A_IWL<11846> A_IWL<11845> A_IWL<11844> A_IWL<11843> A_IWL<11842> A_IWL<11841> A_IWL<11840> A_IWL<11839> A_IWL<11838> A_IWL<11837> A_IWL<11836> A_IWL<11835> A_IWL<11834> A_IWL<11833> A_IWL<11832> A_IWL<11831> A_IWL<11830> A_IWL<11829> A_IWL<11828> A_IWL<11827> A_IWL<11826> A_IWL<11825> A_IWL<11824> A_IWL<11823> A_IWL<11822> A_IWL<11821> A_IWL<11820> A_IWL<11819> A_IWL<11818> A_IWL<11817> A_IWL<11816> A_IWL<11815> A_IWL<11814> A_IWL<11813> A_IWL<11812> A_IWL<11811> A_IWL<11810> A_IWL<11809> A_IWL<11808> A_IWL<11807> A_IWL<11806> A_IWL<11805> A_IWL<11804> A_IWL<11803> A_IWL<11802> A_IWL<11801> A_IWL<11800> A_IWL<11799> A_IWL<11798> A_IWL<11797> A_IWL<11796> A_IWL<11795> A_IWL<11794> A_IWL<11793> A_IWL<11792> A_IWL<11791> A_IWL<11790> A_IWL<11789> A_IWL<11788> A_IWL<11787> A_IWL<11786> A_IWL<11785> A_IWL<11784> A_IWL<11783> A_IWL<11782> A_IWL<11781> A_IWL<11780> A_IWL<11779> A_IWL<11778> A_IWL<11777> A_IWL<11776> A_IWL<12799> A_IWL<12798> A_IWL<12797> A_IWL<12796> A_IWL<12795> A_IWL<12794> A_IWL<12793> A_IWL<12792> A_IWL<12791> A_IWL<12790> A_IWL<12789> A_IWL<12788> A_IWL<12787> A_IWL<12786> A_IWL<12785> A_IWL<12784> A_IWL<12783> A_IWL<12782> A_IWL<12781> A_IWL<12780> A_IWL<12779> A_IWL<12778> A_IWL<12777> A_IWL<12776> A_IWL<12775> A_IWL<12774> A_IWL<12773> A_IWL<12772> A_IWL<12771> A_IWL<12770> A_IWL<12769> A_IWL<12768> A_IWL<12767> A_IWL<12766> A_IWL<12765> A_IWL<12764> A_IWL<12763> A_IWL<12762> A_IWL<12761> A_IWL<12760> A_IWL<12759> A_IWL<12758> A_IWL<12757> A_IWL<12756> A_IWL<12755> A_IWL<12754> A_IWL<12753> A_IWL<12752> A_IWL<12751> A_IWL<12750> A_IWL<12749> A_IWL<12748> A_IWL<12747> A_IWL<12746> A_IWL<12745> A_IWL<12744> A_IWL<12743> A_IWL<12742> A_IWL<12741> A_IWL<12740> A_IWL<12739> A_IWL<12738> A_IWL<12737> A_IWL<12736> A_IWL<12735> A_IWL<12734> A_IWL<12733> A_IWL<12732> A_IWL<12731> A_IWL<12730> A_IWL<12729> A_IWL<12728> A_IWL<12727> A_IWL<12726> A_IWL<12725> A_IWL<12724> A_IWL<12723> A_IWL<12722> A_IWL<12721> A_IWL<12720> A_IWL<12719> A_IWL<12718> A_IWL<12717> A_IWL<12716> A_IWL<12715> A_IWL<12714> A_IWL<12713> A_IWL<12712> A_IWL<12711> A_IWL<12710> A_IWL<12709> A_IWL<12708> A_IWL<12707> A_IWL<12706> A_IWL<12705> A_IWL<12704> A_IWL<12703> A_IWL<12702> A_IWL<12701> A_IWL<12700> A_IWL<12699> A_IWL<12698> A_IWL<12697> A_IWL<12696> A_IWL<12695> A_IWL<12694> A_IWL<12693> A_IWL<12692> A_IWL<12691> A_IWL<12690> A_IWL<12689> A_IWL<12688> A_IWL<12687> A_IWL<12686> A_IWL<12685> A_IWL<12684> A_IWL<12683> A_IWL<12682> A_IWL<12681> A_IWL<12680> A_IWL<12679> A_IWL<12678> A_IWL<12677> A_IWL<12676> A_IWL<12675> A_IWL<12674> A_IWL<12673> A_IWL<12672> A_IWL<12671> A_IWL<12670> A_IWL<12669> A_IWL<12668> A_IWL<12667> A_IWL<12666> A_IWL<12665> A_IWL<12664> A_IWL<12663> A_IWL<12662> A_IWL<12661> A_IWL<12660> A_IWL<12659> A_IWL<12658> A_IWL<12657> A_IWL<12656> A_IWL<12655> A_IWL<12654> A_IWL<12653> A_IWL<12652> A_IWL<12651> A_IWL<12650> A_IWL<12649> A_IWL<12648> A_IWL<12647> A_IWL<12646> A_IWL<12645> A_IWL<12644> A_IWL<12643> A_IWL<12642> A_IWL<12641> A_IWL<12640> A_IWL<12639> A_IWL<12638> A_IWL<12637> A_IWL<12636> A_IWL<12635> A_IWL<12634> A_IWL<12633> A_IWL<12632> A_IWL<12631> A_IWL<12630> A_IWL<12629> A_IWL<12628> A_IWL<12627> A_IWL<12626> A_IWL<12625> A_IWL<12624> A_IWL<12623> A_IWL<12622> A_IWL<12621> A_IWL<12620> A_IWL<12619> A_IWL<12618> A_IWL<12617> A_IWL<12616> A_IWL<12615> A_IWL<12614> A_IWL<12613> A_IWL<12612> A_IWL<12611> A_IWL<12610> A_IWL<12609> A_IWL<12608> A_IWL<12607> A_IWL<12606> A_IWL<12605> A_IWL<12604> A_IWL<12603> A_IWL<12602> A_IWL<12601> A_IWL<12600> A_IWL<12599> A_IWL<12598> A_IWL<12597> A_IWL<12596> A_IWL<12595> A_IWL<12594> A_IWL<12593> A_IWL<12592> A_IWL<12591> A_IWL<12590> A_IWL<12589> A_IWL<12588> A_IWL<12587> A_IWL<12586> A_IWL<12585> A_IWL<12584> A_IWL<12583> A_IWL<12582> A_IWL<12581> A_IWL<12580> A_IWL<12579> A_IWL<12578> A_IWL<12577> A_IWL<12576> A_IWL<12575> A_IWL<12574> A_IWL<12573> A_IWL<12572> A_IWL<12571> A_IWL<12570> A_IWL<12569> A_IWL<12568> A_IWL<12567> A_IWL<12566> A_IWL<12565> A_IWL<12564> A_IWL<12563> A_IWL<12562> A_IWL<12561> A_IWL<12560> A_IWL<12559> A_IWL<12558> A_IWL<12557> A_IWL<12556> A_IWL<12555> A_IWL<12554> A_IWL<12553> A_IWL<12552> A_IWL<12551> A_IWL<12550> A_IWL<12549> A_IWL<12548> A_IWL<12547> A_IWL<12546> A_IWL<12545> A_IWL<12544> A_IWL<12543> A_IWL<12542> A_IWL<12541> A_IWL<12540> A_IWL<12539> A_IWL<12538> A_IWL<12537> A_IWL<12536> A_IWL<12535> A_IWL<12534> A_IWL<12533> A_IWL<12532> A_IWL<12531> A_IWL<12530> A_IWL<12529> A_IWL<12528> A_IWL<12527> A_IWL<12526> A_IWL<12525> A_IWL<12524> A_IWL<12523> A_IWL<12522> A_IWL<12521> A_IWL<12520> A_IWL<12519> A_IWL<12518> A_IWL<12517> A_IWL<12516> A_IWL<12515> A_IWL<12514> A_IWL<12513> A_IWL<12512> A_IWL<12511> A_IWL<12510> A_IWL<12509> A_IWL<12508> A_IWL<12507> A_IWL<12506> A_IWL<12505> A_IWL<12504> A_IWL<12503> A_IWL<12502> A_IWL<12501> A_IWL<12500> A_IWL<12499> A_IWL<12498> A_IWL<12497> A_IWL<12496> A_IWL<12495> A_IWL<12494> A_IWL<12493> A_IWL<12492> A_IWL<12491> A_IWL<12490> A_IWL<12489> A_IWL<12488> A_IWL<12487> A_IWL<12486> A_IWL<12485> A_IWL<12484> A_IWL<12483> A_IWL<12482> A_IWL<12481> A_IWL<12480> A_IWL<12479> A_IWL<12478> A_IWL<12477> A_IWL<12476> A_IWL<12475> A_IWL<12474> A_IWL<12473> A_IWL<12472> A_IWL<12471> A_IWL<12470> A_IWL<12469> A_IWL<12468> A_IWL<12467> A_IWL<12466> A_IWL<12465> A_IWL<12464> A_IWL<12463> A_IWL<12462> A_IWL<12461> A_IWL<12460> A_IWL<12459> A_IWL<12458> A_IWL<12457> A_IWL<12456> A_IWL<12455> A_IWL<12454> A_IWL<12453> A_IWL<12452> A_IWL<12451> A_IWL<12450> A_IWL<12449> A_IWL<12448> A_IWL<12447> A_IWL<12446> A_IWL<12445> A_IWL<12444> A_IWL<12443> A_IWL<12442> A_IWL<12441> A_IWL<12440> A_IWL<12439> A_IWL<12438> A_IWL<12437> A_IWL<12436> A_IWL<12435> A_IWL<12434> A_IWL<12433> A_IWL<12432> A_IWL<12431> A_IWL<12430> A_IWL<12429> A_IWL<12428> A_IWL<12427> A_IWL<12426> A_IWL<12425> A_IWL<12424> A_IWL<12423> A_IWL<12422> A_IWL<12421> A_IWL<12420> A_IWL<12419> A_IWL<12418> A_IWL<12417> A_IWL<12416> A_IWL<12415> A_IWL<12414> A_IWL<12413> A_IWL<12412> A_IWL<12411> A_IWL<12410> A_IWL<12409> A_IWL<12408> A_IWL<12407> A_IWL<12406> A_IWL<12405> A_IWL<12404> A_IWL<12403> A_IWL<12402> A_IWL<12401> A_IWL<12400> A_IWL<12399> A_IWL<12398> A_IWL<12397> A_IWL<12396> A_IWL<12395> A_IWL<12394> A_IWL<12393> A_IWL<12392> A_IWL<12391> A_IWL<12390> A_IWL<12389> A_IWL<12388> A_IWL<12387> A_IWL<12386> A_IWL<12385> A_IWL<12384> A_IWL<12383> A_IWL<12382> A_IWL<12381> A_IWL<12380> A_IWL<12379> A_IWL<12378> A_IWL<12377> A_IWL<12376> A_IWL<12375> A_IWL<12374> A_IWL<12373> A_IWL<12372> A_IWL<12371> A_IWL<12370> A_IWL<12369> A_IWL<12368> A_IWL<12367> A_IWL<12366> A_IWL<12365> A_IWL<12364> A_IWL<12363> A_IWL<12362> A_IWL<12361> A_IWL<12360> A_IWL<12359> A_IWL<12358> A_IWL<12357> A_IWL<12356> A_IWL<12355> A_IWL<12354> A_IWL<12353> A_IWL<12352> A_IWL<12351> A_IWL<12350> A_IWL<12349> A_IWL<12348> A_IWL<12347> A_IWL<12346> A_IWL<12345> A_IWL<12344> A_IWL<12343> A_IWL<12342> A_IWL<12341> A_IWL<12340> A_IWL<12339> A_IWL<12338> A_IWL<12337> A_IWL<12336> A_IWL<12335> A_IWL<12334> A_IWL<12333> A_IWL<12332> A_IWL<12331> A_IWL<12330> A_IWL<12329> A_IWL<12328> A_IWL<12327> A_IWL<12326> A_IWL<12325> A_IWL<12324> A_IWL<12323> A_IWL<12322> A_IWL<12321> A_IWL<12320> A_IWL<12319> A_IWL<12318> A_IWL<12317> A_IWL<12316> A_IWL<12315> A_IWL<12314> A_IWL<12313> A_IWL<12312> A_IWL<12311> A_IWL<12310> A_IWL<12309> A_IWL<12308> A_IWL<12307> A_IWL<12306> A_IWL<12305> A_IWL<12304> A_IWL<12303> A_IWL<12302> A_IWL<12301> A_IWL<12300> A_IWL<12299> A_IWL<12298> A_IWL<12297> A_IWL<12296> A_IWL<12295> A_IWL<12294> A_IWL<12293> A_IWL<12292> A_IWL<12291> A_IWL<12290> A_IWL<12289> A_IWL<12288> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<23> A_BLC<47> A_BLC<46> A_BLC_TOP<47> A_BLC_TOP<46> A_BLT<47> A_BLT<46> A_BLT_TOP<47> A_BLT_TOP<46> A_IWL<11775> A_IWL<11774> A_IWL<11773> A_IWL<11772> A_IWL<11771> A_IWL<11770> A_IWL<11769> A_IWL<11768> A_IWL<11767> A_IWL<11766> A_IWL<11765> A_IWL<11764> A_IWL<11763> A_IWL<11762> A_IWL<11761> A_IWL<11760> A_IWL<11759> A_IWL<11758> A_IWL<11757> A_IWL<11756> A_IWL<11755> A_IWL<11754> A_IWL<11753> A_IWL<11752> A_IWL<11751> A_IWL<11750> A_IWL<11749> A_IWL<11748> A_IWL<11747> A_IWL<11746> A_IWL<11745> A_IWL<11744> A_IWL<11743> A_IWL<11742> A_IWL<11741> A_IWL<11740> A_IWL<11739> A_IWL<11738> A_IWL<11737> A_IWL<11736> A_IWL<11735> A_IWL<11734> A_IWL<11733> A_IWL<11732> A_IWL<11731> A_IWL<11730> A_IWL<11729> A_IWL<11728> A_IWL<11727> A_IWL<11726> A_IWL<11725> A_IWL<11724> A_IWL<11723> A_IWL<11722> A_IWL<11721> A_IWL<11720> A_IWL<11719> A_IWL<11718> A_IWL<11717> A_IWL<11716> A_IWL<11715> A_IWL<11714> A_IWL<11713> A_IWL<11712> A_IWL<11711> A_IWL<11710> A_IWL<11709> A_IWL<11708> A_IWL<11707> A_IWL<11706> A_IWL<11705> A_IWL<11704> A_IWL<11703> A_IWL<11702> A_IWL<11701> A_IWL<11700> A_IWL<11699> A_IWL<11698> A_IWL<11697> A_IWL<11696> A_IWL<11695> A_IWL<11694> A_IWL<11693> A_IWL<11692> A_IWL<11691> A_IWL<11690> A_IWL<11689> A_IWL<11688> A_IWL<11687> A_IWL<11686> A_IWL<11685> A_IWL<11684> A_IWL<11683> A_IWL<11682> A_IWL<11681> A_IWL<11680> A_IWL<11679> A_IWL<11678> A_IWL<11677> A_IWL<11676> A_IWL<11675> A_IWL<11674> A_IWL<11673> A_IWL<11672> A_IWL<11671> A_IWL<11670> A_IWL<11669> A_IWL<11668> A_IWL<11667> A_IWL<11666> A_IWL<11665> A_IWL<11664> A_IWL<11663> A_IWL<11662> A_IWL<11661> A_IWL<11660> A_IWL<11659> A_IWL<11658> A_IWL<11657> A_IWL<11656> A_IWL<11655> A_IWL<11654> A_IWL<11653> A_IWL<11652> A_IWL<11651> A_IWL<11650> A_IWL<11649> A_IWL<11648> A_IWL<11647> A_IWL<11646> A_IWL<11645> A_IWL<11644> A_IWL<11643> A_IWL<11642> A_IWL<11641> A_IWL<11640> A_IWL<11639> A_IWL<11638> A_IWL<11637> A_IWL<11636> A_IWL<11635> A_IWL<11634> A_IWL<11633> A_IWL<11632> A_IWL<11631> A_IWL<11630> A_IWL<11629> A_IWL<11628> A_IWL<11627> A_IWL<11626> A_IWL<11625> A_IWL<11624> A_IWL<11623> A_IWL<11622> A_IWL<11621> A_IWL<11620> A_IWL<11619> A_IWL<11618> A_IWL<11617> A_IWL<11616> A_IWL<11615> A_IWL<11614> A_IWL<11613> A_IWL<11612> A_IWL<11611> A_IWL<11610> A_IWL<11609> A_IWL<11608> A_IWL<11607> A_IWL<11606> A_IWL<11605> A_IWL<11604> A_IWL<11603> A_IWL<11602> A_IWL<11601> A_IWL<11600> A_IWL<11599> A_IWL<11598> A_IWL<11597> A_IWL<11596> A_IWL<11595> A_IWL<11594> A_IWL<11593> A_IWL<11592> A_IWL<11591> A_IWL<11590> A_IWL<11589> A_IWL<11588> A_IWL<11587> A_IWL<11586> A_IWL<11585> A_IWL<11584> A_IWL<11583> A_IWL<11582> A_IWL<11581> A_IWL<11580> A_IWL<11579> A_IWL<11578> A_IWL<11577> A_IWL<11576> A_IWL<11575> A_IWL<11574> A_IWL<11573> A_IWL<11572> A_IWL<11571> A_IWL<11570> A_IWL<11569> A_IWL<11568> A_IWL<11567> A_IWL<11566> A_IWL<11565> A_IWL<11564> A_IWL<11563> A_IWL<11562> A_IWL<11561> A_IWL<11560> A_IWL<11559> A_IWL<11558> A_IWL<11557> A_IWL<11556> A_IWL<11555> A_IWL<11554> A_IWL<11553> A_IWL<11552> A_IWL<11551> A_IWL<11550> A_IWL<11549> A_IWL<11548> A_IWL<11547> A_IWL<11546> A_IWL<11545> A_IWL<11544> A_IWL<11543> A_IWL<11542> A_IWL<11541> A_IWL<11540> A_IWL<11539> A_IWL<11538> A_IWL<11537> A_IWL<11536> A_IWL<11535> A_IWL<11534> A_IWL<11533> A_IWL<11532> A_IWL<11531> A_IWL<11530> A_IWL<11529> A_IWL<11528> A_IWL<11527> A_IWL<11526> A_IWL<11525> A_IWL<11524> A_IWL<11523> A_IWL<11522> A_IWL<11521> A_IWL<11520> A_IWL<11519> A_IWL<11518> A_IWL<11517> A_IWL<11516> A_IWL<11515> A_IWL<11514> A_IWL<11513> A_IWL<11512> A_IWL<11511> A_IWL<11510> A_IWL<11509> A_IWL<11508> A_IWL<11507> A_IWL<11506> A_IWL<11505> A_IWL<11504> A_IWL<11503> A_IWL<11502> A_IWL<11501> A_IWL<11500> A_IWL<11499> A_IWL<11498> A_IWL<11497> A_IWL<11496> A_IWL<11495> A_IWL<11494> A_IWL<11493> A_IWL<11492> A_IWL<11491> A_IWL<11490> A_IWL<11489> A_IWL<11488> A_IWL<11487> A_IWL<11486> A_IWL<11485> A_IWL<11484> A_IWL<11483> A_IWL<11482> A_IWL<11481> A_IWL<11480> A_IWL<11479> A_IWL<11478> A_IWL<11477> A_IWL<11476> A_IWL<11475> A_IWL<11474> A_IWL<11473> A_IWL<11472> A_IWL<11471> A_IWL<11470> A_IWL<11469> A_IWL<11468> A_IWL<11467> A_IWL<11466> A_IWL<11465> A_IWL<11464> A_IWL<11463> A_IWL<11462> A_IWL<11461> A_IWL<11460> A_IWL<11459> A_IWL<11458> A_IWL<11457> A_IWL<11456> A_IWL<11455> A_IWL<11454> A_IWL<11453> A_IWL<11452> A_IWL<11451> A_IWL<11450> A_IWL<11449> A_IWL<11448> A_IWL<11447> A_IWL<11446> A_IWL<11445> A_IWL<11444> A_IWL<11443> A_IWL<11442> A_IWL<11441> A_IWL<11440> A_IWL<11439> A_IWL<11438> A_IWL<11437> A_IWL<11436> A_IWL<11435> A_IWL<11434> A_IWL<11433> A_IWL<11432> A_IWL<11431> A_IWL<11430> A_IWL<11429> A_IWL<11428> A_IWL<11427> A_IWL<11426> A_IWL<11425> A_IWL<11424> A_IWL<11423> A_IWL<11422> A_IWL<11421> A_IWL<11420> A_IWL<11419> A_IWL<11418> A_IWL<11417> A_IWL<11416> A_IWL<11415> A_IWL<11414> A_IWL<11413> A_IWL<11412> A_IWL<11411> A_IWL<11410> A_IWL<11409> A_IWL<11408> A_IWL<11407> A_IWL<11406> A_IWL<11405> A_IWL<11404> A_IWL<11403> A_IWL<11402> A_IWL<11401> A_IWL<11400> A_IWL<11399> A_IWL<11398> A_IWL<11397> A_IWL<11396> A_IWL<11395> A_IWL<11394> A_IWL<11393> A_IWL<11392> A_IWL<11391> A_IWL<11390> A_IWL<11389> A_IWL<11388> A_IWL<11387> A_IWL<11386> A_IWL<11385> A_IWL<11384> A_IWL<11383> A_IWL<11382> A_IWL<11381> A_IWL<11380> A_IWL<11379> A_IWL<11378> A_IWL<11377> A_IWL<11376> A_IWL<11375> A_IWL<11374> A_IWL<11373> A_IWL<11372> A_IWL<11371> A_IWL<11370> A_IWL<11369> A_IWL<11368> A_IWL<11367> A_IWL<11366> A_IWL<11365> A_IWL<11364> A_IWL<11363> A_IWL<11362> A_IWL<11361> A_IWL<11360> A_IWL<11359> A_IWL<11358> A_IWL<11357> A_IWL<11356> A_IWL<11355> A_IWL<11354> A_IWL<11353> A_IWL<11352> A_IWL<11351> A_IWL<11350> A_IWL<11349> A_IWL<11348> A_IWL<11347> A_IWL<11346> A_IWL<11345> A_IWL<11344> A_IWL<11343> A_IWL<11342> A_IWL<11341> A_IWL<11340> A_IWL<11339> A_IWL<11338> A_IWL<11337> A_IWL<11336> A_IWL<11335> A_IWL<11334> A_IWL<11333> A_IWL<11332> A_IWL<11331> A_IWL<11330> A_IWL<11329> A_IWL<11328> A_IWL<11327> A_IWL<11326> A_IWL<11325> A_IWL<11324> A_IWL<11323> A_IWL<11322> A_IWL<11321> A_IWL<11320> A_IWL<11319> A_IWL<11318> A_IWL<11317> A_IWL<11316> A_IWL<11315> A_IWL<11314> A_IWL<11313> A_IWL<11312> A_IWL<11311> A_IWL<11310> A_IWL<11309> A_IWL<11308> A_IWL<11307> A_IWL<11306> A_IWL<11305> A_IWL<11304> A_IWL<11303> A_IWL<11302> A_IWL<11301> A_IWL<11300> A_IWL<11299> A_IWL<11298> A_IWL<11297> A_IWL<11296> A_IWL<11295> A_IWL<11294> A_IWL<11293> A_IWL<11292> A_IWL<11291> A_IWL<11290> A_IWL<11289> A_IWL<11288> A_IWL<11287> A_IWL<11286> A_IWL<11285> A_IWL<11284> A_IWL<11283> A_IWL<11282> A_IWL<11281> A_IWL<11280> A_IWL<11279> A_IWL<11278> A_IWL<11277> A_IWL<11276> A_IWL<11275> A_IWL<11274> A_IWL<11273> A_IWL<11272> A_IWL<11271> A_IWL<11270> A_IWL<11269> A_IWL<11268> A_IWL<11267> A_IWL<11266> A_IWL<11265> A_IWL<11264> A_IWL<12287> A_IWL<12286> A_IWL<12285> A_IWL<12284> A_IWL<12283> A_IWL<12282> A_IWL<12281> A_IWL<12280> A_IWL<12279> A_IWL<12278> A_IWL<12277> A_IWL<12276> A_IWL<12275> A_IWL<12274> A_IWL<12273> A_IWL<12272> A_IWL<12271> A_IWL<12270> A_IWL<12269> A_IWL<12268> A_IWL<12267> A_IWL<12266> A_IWL<12265> A_IWL<12264> A_IWL<12263> A_IWL<12262> A_IWL<12261> A_IWL<12260> A_IWL<12259> A_IWL<12258> A_IWL<12257> A_IWL<12256> A_IWL<12255> A_IWL<12254> A_IWL<12253> A_IWL<12252> A_IWL<12251> A_IWL<12250> A_IWL<12249> A_IWL<12248> A_IWL<12247> A_IWL<12246> A_IWL<12245> A_IWL<12244> A_IWL<12243> A_IWL<12242> A_IWL<12241> A_IWL<12240> A_IWL<12239> A_IWL<12238> A_IWL<12237> A_IWL<12236> A_IWL<12235> A_IWL<12234> A_IWL<12233> A_IWL<12232> A_IWL<12231> A_IWL<12230> A_IWL<12229> A_IWL<12228> A_IWL<12227> A_IWL<12226> A_IWL<12225> A_IWL<12224> A_IWL<12223> A_IWL<12222> A_IWL<12221> A_IWL<12220> A_IWL<12219> A_IWL<12218> A_IWL<12217> A_IWL<12216> A_IWL<12215> A_IWL<12214> A_IWL<12213> A_IWL<12212> A_IWL<12211> A_IWL<12210> A_IWL<12209> A_IWL<12208> A_IWL<12207> A_IWL<12206> A_IWL<12205> A_IWL<12204> A_IWL<12203> A_IWL<12202> A_IWL<12201> A_IWL<12200> A_IWL<12199> A_IWL<12198> A_IWL<12197> A_IWL<12196> A_IWL<12195> A_IWL<12194> A_IWL<12193> A_IWL<12192> A_IWL<12191> A_IWL<12190> A_IWL<12189> A_IWL<12188> A_IWL<12187> A_IWL<12186> A_IWL<12185> A_IWL<12184> A_IWL<12183> A_IWL<12182> A_IWL<12181> A_IWL<12180> A_IWL<12179> A_IWL<12178> A_IWL<12177> A_IWL<12176> A_IWL<12175> A_IWL<12174> A_IWL<12173> A_IWL<12172> A_IWL<12171> A_IWL<12170> A_IWL<12169> A_IWL<12168> A_IWL<12167> A_IWL<12166> A_IWL<12165> A_IWL<12164> A_IWL<12163> A_IWL<12162> A_IWL<12161> A_IWL<12160> A_IWL<12159> A_IWL<12158> A_IWL<12157> A_IWL<12156> A_IWL<12155> A_IWL<12154> A_IWL<12153> A_IWL<12152> A_IWL<12151> A_IWL<12150> A_IWL<12149> A_IWL<12148> A_IWL<12147> A_IWL<12146> A_IWL<12145> A_IWL<12144> A_IWL<12143> A_IWL<12142> A_IWL<12141> A_IWL<12140> A_IWL<12139> A_IWL<12138> A_IWL<12137> A_IWL<12136> A_IWL<12135> A_IWL<12134> A_IWL<12133> A_IWL<12132> A_IWL<12131> A_IWL<12130> A_IWL<12129> A_IWL<12128> A_IWL<12127> A_IWL<12126> A_IWL<12125> A_IWL<12124> A_IWL<12123> A_IWL<12122> A_IWL<12121> A_IWL<12120> A_IWL<12119> A_IWL<12118> A_IWL<12117> A_IWL<12116> A_IWL<12115> A_IWL<12114> A_IWL<12113> A_IWL<12112> A_IWL<12111> A_IWL<12110> A_IWL<12109> A_IWL<12108> A_IWL<12107> A_IWL<12106> A_IWL<12105> A_IWL<12104> A_IWL<12103> A_IWL<12102> A_IWL<12101> A_IWL<12100> A_IWL<12099> A_IWL<12098> A_IWL<12097> A_IWL<12096> A_IWL<12095> A_IWL<12094> A_IWL<12093> A_IWL<12092> A_IWL<12091> A_IWL<12090> A_IWL<12089> A_IWL<12088> A_IWL<12087> A_IWL<12086> A_IWL<12085> A_IWL<12084> A_IWL<12083> A_IWL<12082> A_IWL<12081> A_IWL<12080> A_IWL<12079> A_IWL<12078> A_IWL<12077> A_IWL<12076> A_IWL<12075> A_IWL<12074> A_IWL<12073> A_IWL<12072> A_IWL<12071> A_IWL<12070> A_IWL<12069> A_IWL<12068> A_IWL<12067> A_IWL<12066> A_IWL<12065> A_IWL<12064> A_IWL<12063> A_IWL<12062> A_IWL<12061> A_IWL<12060> A_IWL<12059> A_IWL<12058> A_IWL<12057> A_IWL<12056> A_IWL<12055> A_IWL<12054> A_IWL<12053> A_IWL<12052> A_IWL<12051> A_IWL<12050> A_IWL<12049> A_IWL<12048> A_IWL<12047> A_IWL<12046> A_IWL<12045> A_IWL<12044> A_IWL<12043> A_IWL<12042> A_IWL<12041> A_IWL<12040> A_IWL<12039> A_IWL<12038> A_IWL<12037> A_IWL<12036> A_IWL<12035> A_IWL<12034> A_IWL<12033> A_IWL<12032> A_IWL<12031> A_IWL<12030> A_IWL<12029> A_IWL<12028> A_IWL<12027> A_IWL<12026> A_IWL<12025> A_IWL<12024> A_IWL<12023> A_IWL<12022> A_IWL<12021> A_IWL<12020> A_IWL<12019> A_IWL<12018> A_IWL<12017> A_IWL<12016> A_IWL<12015> A_IWL<12014> A_IWL<12013> A_IWL<12012> A_IWL<12011> A_IWL<12010> A_IWL<12009> A_IWL<12008> A_IWL<12007> A_IWL<12006> A_IWL<12005> A_IWL<12004> A_IWL<12003> A_IWL<12002> A_IWL<12001> A_IWL<12000> A_IWL<11999> A_IWL<11998> A_IWL<11997> A_IWL<11996> A_IWL<11995> A_IWL<11994> A_IWL<11993> A_IWL<11992> A_IWL<11991> A_IWL<11990> A_IWL<11989> A_IWL<11988> A_IWL<11987> A_IWL<11986> A_IWL<11985> A_IWL<11984> A_IWL<11983> A_IWL<11982> A_IWL<11981> A_IWL<11980> A_IWL<11979> A_IWL<11978> A_IWL<11977> A_IWL<11976> A_IWL<11975> A_IWL<11974> A_IWL<11973> A_IWL<11972> A_IWL<11971> A_IWL<11970> A_IWL<11969> A_IWL<11968> A_IWL<11967> A_IWL<11966> A_IWL<11965> A_IWL<11964> A_IWL<11963> A_IWL<11962> A_IWL<11961> A_IWL<11960> A_IWL<11959> A_IWL<11958> A_IWL<11957> A_IWL<11956> A_IWL<11955> A_IWL<11954> A_IWL<11953> A_IWL<11952> A_IWL<11951> A_IWL<11950> A_IWL<11949> A_IWL<11948> A_IWL<11947> A_IWL<11946> A_IWL<11945> A_IWL<11944> A_IWL<11943> A_IWL<11942> A_IWL<11941> A_IWL<11940> A_IWL<11939> A_IWL<11938> A_IWL<11937> A_IWL<11936> A_IWL<11935> A_IWL<11934> A_IWL<11933> A_IWL<11932> A_IWL<11931> A_IWL<11930> A_IWL<11929> A_IWL<11928> A_IWL<11927> A_IWL<11926> A_IWL<11925> A_IWL<11924> A_IWL<11923> A_IWL<11922> A_IWL<11921> A_IWL<11920> A_IWL<11919> A_IWL<11918> A_IWL<11917> A_IWL<11916> A_IWL<11915> A_IWL<11914> A_IWL<11913> A_IWL<11912> A_IWL<11911> A_IWL<11910> A_IWL<11909> A_IWL<11908> A_IWL<11907> A_IWL<11906> A_IWL<11905> A_IWL<11904> A_IWL<11903> A_IWL<11902> A_IWL<11901> A_IWL<11900> A_IWL<11899> A_IWL<11898> A_IWL<11897> A_IWL<11896> A_IWL<11895> A_IWL<11894> A_IWL<11893> A_IWL<11892> A_IWL<11891> A_IWL<11890> A_IWL<11889> A_IWL<11888> A_IWL<11887> A_IWL<11886> A_IWL<11885> A_IWL<11884> A_IWL<11883> A_IWL<11882> A_IWL<11881> A_IWL<11880> A_IWL<11879> A_IWL<11878> A_IWL<11877> A_IWL<11876> A_IWL<11875> A_IWL<11874> A_IWL<11873> A_IWL<11872> A_IWL<11871> A_IWL<11870> A_IWL<11869> A_IWL<11868> A_IWL<11867> A_IWL<11866> A_IWL<11865> A_IWL<11864> A_IWL<11863> A_IWL<11862> A_IWL<11861> A_IWL<11860> A_IWL<11859> A_IWL<11858> A_IWL<11857> A_IWL<11856> A_IWL<11855> A_IWL<11854> A_IWL<11853> A_IWL<11852> A_IWL<11851> A_IWL<11850> A_IWL<11849> A_IWL<11848> A_IWL<11847> A_IWL<11846> A_IWL<11845> A_IWL<11844> A_IWL<11843> A_IWL<11842> A_IWL<11841> A_IWL<11840> A_IWL<11839> A_IWL<11838> A_IWL<11837> A_IWL<11836> A_IWL<11835> A_IWL<11834> A_IWL<11833> A_IWL<11832> A_IWL<11831> A_IWL<11830> A_IWL<11829> A_IWL<11828> A_IWL<11827> A_IWL<11826> A_IWL<11825> A_IWL<11824> A_IWL<11823> A_IWL<11822> A_IWL<11821> A_IWL<11820> A_IWL<11819> A_IWL<11818> A_IWL<11817> A_IWL<11816> A_IWL<11815> A_IWL<11814> A_IWL<11813> A_IWL<11812> A_IWL<11811> A_IWL<11810> A_IWL<11809> A_IWL<11808> A_IWL<11807> A_IWL<11806> A_IWL<11805> A_IWL<11804> A_IWL<11803> A_IWL<11802> A_IWL<11801> A_IWL<11800> A_IWL<11799> A_IWL<11798> A_IWL<11797> A_IWL<11796> A_IWL<11795> A_IWL<11794> A_IWL<11793> A_IWL<11792> A_IWL<11791> A_IWL<11790> A_IWL<11789> A_IWL<11788> A_IWL<11787> A_IWL<11786> A_IWL<11785> A_IWL<11784> A_IWL<11783> A_IWL<11782> A_IWL<11781> A_IWL<11780> A_IWL<11779> A_IWL<11778> A_IWL<11777> A_IWL<11776> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<22> A_BLC<45> A_BLC<44> A_BLC_TOP<45> A_BLC_TOP<44> A_BLT<45> A_BLT<44> A_BLT_TOP<45> A_BLT_TOP<44> A_IWL<11263> A_IWL<11262> A_IWL<11261> A_IWL<11260> A_IWL<11259> A_IWL<11258> A_IWL<11257> A_IWL<11256> A_IWL<11255> A_IWL<11254> A_IWL<11253> A_IWL<11252> A_IWL<11251> A_IWL<11250> A_IWL<11249> A_IWL<11248> A_IWL<11247> A_IWL<11246> A_IWL<11245> A_IWL<11244> A_IWL<11243> A_IWL<11242> A_IWL<11241> A_IWL<11240> A_IWL<11239> A_IWL<11238> A_IWL<11237> A_IWL<11236> A_IWL<11235> A_IWL<11234> A_IWL<11233> A_IWL<11232> A_IWL<11231> A_IWL<11230> A_IWL<11229> A_IWL<11228> A_IWL<11227> A_IWL<11226> A_IWL<11225> A_IWL<11224> A_IWL<11223> A_IWL<11222> A_IWL<11221> A_IWL<11220> A_IWL<11219> A_IWL<11218> A_IWL<11217> A_IWL<11216> A_IWL<11215> A_IWL<11214> A_IWL<11213> A_IWL<11212> A_IWL<11211> A_IWL<11210> A_IWL<11209> A_IWL<11208> A_IWL<11207> A_IWL<11206> A_IWL<11205> A_IWL<11204> A_IWL<11203> A_IWL<11202> A_IWL<11201> A_IWL<11200> A_IWL<11199> A_IWL<11198> A_IWL<11197> A_IWL<11196> A_IWL<11195> A_IWL<11194> A_IWL<11193> A_IWL<11192> A_IWL<11191> A_IWL<11190> A_IWL<11189> A_IWL<11188> A_IWL<11187> A_IWL<11186> A_IWL<11185> A_IWL<11184> A_IWL<11183> A_IWL<11182> A_IWL<11181> A_IWL<11180> A_IWL<11179> A_IWL<11178> A_IWL<11177> A_IWL<11176> A_IWL<11175> A_IWL<11174> A_IWL<11173> A_IWL<11172> A_IWL<11171> A_IWL<11170> A_IWL<11169> A_IWL<11168> A_IWL<11167> A_IWL<11166> A_IWL<11165> A_IWL<11164> A_IWL<11163> A_IWL<11162> A_IWL<11161> A_IWL<11160> A_IWL<11159> A_IWL<11158> A_IWL<11157> A_IWL<11156> A_IWL<11155> A_IWL<11154> A_IWL<11153> A_IWL<11152> A_IWL<11151> A_IWL<11150> A_IWL<11149> A_IWL<11148> A_IWL<11147> A_IWL<11146> A_IWL<11145> A_IWL<11144> A_IWL<11143> A_IWL<11142> A_IWL<11141> A_IWL<11140> A_IWL<11139> A_IWL<11138> A_IWL<11137> A_IWL<11136> A_IWL<11135> A_IWL<11134> A_IWL<11133> A_IWL<11132> A_IWL<11131> A_IWL<11130> A_IWL<11129> A_IWL<11128> A_IWL<11127> A_IWL<11126> A_IWL<11125> A_IWL<11124> A_IWL<11123> A_IWL<11122> A_IWL<11121> A_IWL<11120> A_IWL<11119> A_IWL<11118> A_IWL<11117> A_IWL<11116> A_IWL<11115> A_IWL<11114> A_IWL<11113> A_IWL<11112> A_IWL<11111> A_IWL<11110> A_IWL<11109> A_IWL<11108> A_IWL<11107> A_IWL<11106> A_IWL<11105> A_IWL<11104> A_IWL<11103> A_IWL<11102> A_IWL<11101> A_IWL<11100> A_IWL<11099> A_IWL<11098> A_IWL<11097> A_IWL<11096> A_IWL<11095> A_IWL<11094> A_IWL<11093> A_IWL<11092> A_IWL<11091> A_IWL<11090> A_IWL<11089> A_IWL<11088> A_IWL<11087> A_IWL<11086> A_IWL<11085> A_IWL<11084> A_IWL<11083> A_IWL<11082> A_IWL<11081> A_IWL<11080> A_IWL<11079> A_IWL<11078> A_IWL<11077> A_IWL<11076> A_IWL<11075> A_IWL<11074> A_IWL<11073> A_IWL<11072> A_IWL<11071> A_IWL<11070> A_IWL<11069> A_IWL<11068> A_IWL<11067> A_IWL<11066> A_IWL<11065> A_IWL<11064> A_IWL<11063> A_IWL<11062> A_IWL<11061> A_IWL<11060> A_IWL<11059> A_IWL<11058> A_IWL<11057> A_IWL<11056> A_IWL<11055> A_IWL<11054> A_IWL<11053> A_IWL<11052> A_IWL<11051> A_IWL<11050> A_IWL<11049> A_IWL<11048> A_IWL<11047> A_IWL<11046> A_IWL<11045> A_IWL<11044> A_IWL<11043> A_IWL<11042> A_IWL<11041> A_IWL<11040> A_IWL<11039> A_IWL<11038> A_IWL<11037> A_IWL<11036> A_IWL<11035> A_IWL<11034> A_IWL<11033> A_IWL<11032> A_IWL<11031> A_IWL<11030> A_IWL<11029> A_IWL<11028> A_IWL<11027> A_IWL<11026> A_IWL<11025> A_IWL<11024> A_IWL<11023> A_IWL<11022> A_IWL<11021> A_IWL<11020> A_IWL<11019> A_IWL<11018> A_IWL<11017> A_IWL<11016> A_IWL<11015> A_IWL<11014> A_IWL<11013> A_IWL<11012> A_IWL<11011> A_IWL<11010> A_IWL<11009> A_IWL<11008> A_IWL<11007> A_IWL<11006> A_IWL<11005> A_IWL<11004> A_IWL<11003> A_IWL<11002> A_IWL<11001> A_IWL<11000> A_IWL<10999> A_IWL<10998> A_IWL<10997> A_IWL<10996> A_IWL<10995> A_IWL<10994> A_IWL<10993> A_IWL<10992> A_IWL<10991> A_IWL<10990> A_IWL<10989> A_IWL<10988> A_IWL<10987> A_IWL<10986> A_IWL<10985> A_IWL<10984> A_IWL<10983> A_IWL<10982> A_IWL<10981> A_IWL<10980> A_IWL<10979> A_IWL<10978> A_IWL<10977> A_IWL<10976> A_IWL<10975> A_IWL<10974> A_IWL<10973> A_IWL<10972> A_IWL<10971> A_IWL<10970> A_IWL<10969> A_IWL<10968> A_IWL<10967> A_IWL<10966> A_IWL<10965> A_IWL<10964> A_IWL<10963> A_IWL<10962> A_IWL<10961> A_IWL<10960> A_IWL<10959> A_IWL<10958> A_IWL<10957> A_IWL<10956> A_IWL<10955> A_IWL<10954> A_IWL<10953> A_IWL<10952> A_IWL<10951> A_IWL<10950> A_IWL<10949> A_IWL<10948> A_IWL<10947> A_IWL<10946> A_IWL<10945> A_IWL<10944> A_IWL<10943> A_IWL<10942> A_IWL<10941> A_IWL<10940> A_IWL<10939> A_IWL<10938> A_IWL<10937> A_IWL<10936> A_IWL<10935> A_IWL<10934> A_IWL<10933> A_IWL<10932> A_IWL<10931> A_IWL<10930> A_IWL<10929> A_IWL<10928> A_IWL<10927> A_IWL<10926> A_IWL<10925> A_IWL<10924> A_IWL<10923> A_IWL<10922> A_IWL<10921> A_IWL<10920> A_IWL<10919> A_IWL<10918> A_IWL<10917> A_IWL<10916> A_IWL<10915> A_IWL<10914> A_IWL<10913> A_IWL<10912> A_IWL<10911> A_IWL<10910> A_IWL<10909> A_IWL<10908> A_IWL<10907> A_IWL<10906> A_IWL<10905> A_IWL<10904> A_IWL<10903> A_IWL<10902> A_IWL<10901> A_IWL<10900> A_IWL<10899> A_IWL<10898> A_IWL<10897> A_IWL<10896> A_IWL<10895> A_IWL<10894> A_IWL<10893> A_IWL<10892> A_IWL<10891> A_IWL<10890> A_IWL<10889> A_IWL<10888> A_IWL<10887> A_IWL<10886> A_IWL<10885> A_IWL<10884> A_IWL<10883> A_IWL<10882> A_IWL<10881> A_IWL<10880> A_IWL<10879> A_IWL<10878> A_IWL<10877> A_IWL<10876> A_IWL<10875> A_IWL<10874> A_IWL<10873> A_IWL<10872> A_IWL<10871> A_IWL<10870> A_IWL<10869> A_IWL<10868> A_IWL<10867> A_IWL<10866> A_IWL<10865> A_IWL<10864> A_IWL<10863> A_IWL<10862> A_IWL<10861> A_IWL<10860> A_IWL<10859> A_IWL<10858> A_IWL<10857> A_IWL<10856> A_IWL<10855> A_IWL<10854> A_IWL<10853> A_IWL<10852> A_IWL<10851> A_IWL<10850> A_IWL<10849> A_IWL<10848> A_IWL<10847> A_IWL<10846> A_IWL<10845> A_IWL<10844> A_IWL<10843> A_IWL<10842> A_IWL<10841> A_IWL<10840> A_IWL<10839> A_IWL<10838> A_IWL<10837> A_IWL<10836> A_IWL<10835> A_IWL<10834> A_IWL<10833> A_IWL<10832> A_IWL<10831> A_IWL<10830> A_IWL<10829> A_IWL<10828> A_IWL<10827> A_IWL<10826> A_IWL<10825> A_IWL<10824> A_IWL<10823> A_IWL<10822> A_IWL<10821> A_IWL<10820> A_IWL<10819> A_IWL<10818> A_IWL<10817> A_IWL<10816> A_IWL<10815> A_IWL<10814> A_IWL<10813> A_IWL<10812> A_IWL<10811> A_IWL<10810> A_IWL<10809> A_IWL<10808> A_IWL<10807> A_IWL<10806> A_IWL<10805> A_IWL<10804> A_IWL<10803> A_IWL<10802> A_IWL<10801> A_IWL<10800> A_IWL<10799> A_IWL<10798> A_IWL<10797> A_IWL<10796> A_IWL<10795> A_IWL<10794> A_IWL<10793> A_IWL<10792> A_IWL<10791> A_IWL<10790> A_IWL<10789> A_IWL<10788> A_IWL<10787> A_IWL<10786> A_IWL<10785> A_IWL<10784> A_IWL<10783> A_IWL<10782> A_IWL<10781> A_IWL<10780> A_IWL<10779> A_IWL<10778> A_IWL<10777> A_IWL<10776> A_IWL<10775> A_IWL<10774> A_IWL<10773> A_IWL<10772> A_IWL<10771> A_IWL<10770> A_IWL<10769> A_IWL<10768> A_IWL<10767> A_IWL<10766> A_IWL<10765> A_IWL<10764> A_IWL<10763> A_IWL<10762> A_IWL<10761> A_IWL<10760> A_IWL<10759> A_IWL<10758> A_IWL<10757> A_IWL<10756> A_IWL<10755> A_IWL<10754> A_IWL<10753> A_IWL<10752> A_IWL<11775> A_IWL<11774> A_IWL<11773> A_IWL<11772> A_IWL<11771> A_IWL<11770> A_IWL<11769> A_IWL<11768> A_IWL<11767> A_IWL<11766> A_IWL<11765> A_IWL<11764> A_IWL<11763> A_IWL<11762> A_IWL<11761> A_IWL<11760> A_IWL<11759> A_IWL<11758> A_IWL<11757> A_IWL<11756> A_IWL<11755> A_IWL<11754> A_IWL<11753> A_IWL<11752> A_IWL<11751> A_IWL<11750> A_IWL<11749> A_IWL<11748> A_IWL<11747> A_IWL<11746> A_IWL<11745> A_IWL<11744> A_IWL<11743> A_IWL<11742> A_IWL<11741> A_IWL<11740> A_IWL<11739> A_IWL<11738> A_IWL<11737> A_IWL<11736> A_IWL<11735> A_IWL<11734> A_IWL<11733> A_IWL<11732> A_IWL<11731> A_IWL<11730> A_IWL<11729> A_IWL<11728> A_IWL<11727> A_IWL<11726> A_IWL<11725> A_IWL<11724> A_IWL<11723> A_IWL<11722> A_IWL<11721> A_IWL<11720> A_IWL<11719> A_IWL<11718> A_IWL<11717> A_IWL<11716> A_IWL<11715> A_IWL<11714> A_IWL<11713> A_IWL<11712> A_IWL<11711> A_IWL<11710> A_IWL<11709> A_IWL<11708> A_IWL<11707> A_IWL<11706> A_IWL<11705> A_IWL<11704> A_IWL<11703> A_IWL<11702> A_IWL<11701> A_IWL<11700> A_IWL<11699> A_IWL<11698> A_IWL<11697> A_IWL<11696> A_IWL<11695> A_IWL<11694> A_IWL<11693> A_IWL<11692> A_IWL<11691> A_IWL<11690> A_IWL<11689> A_IWL<11688> A_IWL<11687> A_IWL<11686> A_IWL<11685> A_IWL<11684> A_IWL<11683> A_IWL<11682> A_IWL<11681> A_IWL<11680> A_IWL<11679> A_IWL<11678> A_IWL<11677> A_IWL<11676> A_IWL<11675> A_IWL<11674> A_IWL<11673> A_IWL<11672> A_IWL<11671> A_IWL<11670> A_IWL<11669> A_IWL<11668> A_IWL<11667> A_IWL<11666> A_IWL<11665> A_IWL<11664> A_IWL<11663> A_IWL<11662> A_IWL<11661> A_IWL<11660> A_IWL<11659> A_IWL<11658> A_IWL<11657> A_IWL<11656> A_IWL<11655> A_IWL<11654> A_IWL<11653> A_IWL<11652> A_IWL<11651> A_IWL<11650> A_IWL<11649> A_IWL<11648> A_IWL<11647> A_IWL<11646> A_IWL<11645> A_IWL<11644> A_IWL<11643> A_IWL<11642> A_IWL<11641> A_IWL<11640> A_IWL<11639> A_IWL<11638> A_IWL<11637> A_IWL<11636> A_IWL<11635> A_IWL<11634> A_IWL<11633> A_IWL<11632> A_IWL<11631> A_IWL<11630> A_IWL<11629> A_IWL<11628> A_IWL<11627> A_IWL<11626> A_IWL<11625> A_IWL<11624> A_IWL<11623> A_IWL<11622> A_IWL<11621> A_IWL<11620> A_IWL<11619> A_IWL<11618> A_IWL<11617> A_IWL<11616> A_IWL<11615> A_IWL<11614> A_IWL<11613> A_IWL<11612> A_IWL<11611> A_IWL<11610> A_IWL<11609> A_IWL<11608> A_IWL<11607> A_IWL<11606> A_IWL<11605> A_IWL<11604> A_IWL<11603> A_IWL<11602> A_IWL<11601> A_IWL<11600> A_IWL<11599> A_IWL<11598> A_IWL<11597> A_IWL<11596> A_IWL<11595> A_IWL<11594> A_IWL<11593> A_IWL<11592> A_IWL<11591> A_IWL<11590> A_IWL<11589> A_IWL<11588> A_IWL<11587> A_IWL<11586> A_IWL<11585> A_IWL<11584> A_IWL<11583> A_IWL<11582> A_IWL<11581> A_IWL<11580> A_IWL<11579> A_IWL<11578> A_IWL<11577> A_IWL<11576> A_IWL<11575> A_IWL<11574> A_IWL<11573> A_IWL<11572> A_IWL<11571> A_IWL<11570> A_IWL<11569> A_IWL<11568> A_IWL<11567> A_IWL<11566> A_IWL<11565> A_IWL<11564> A_IWL<11563> A_IWL<11562> A_IWL<11561> A_IWL<11560> A_IWL<11559> A_IWL<11558> A_IWL<11557> A_IWL<11556> A_IWL<11555> A_IWL<11554> A_IWL<11553> A_IWL<11552> A_IWL<11551> A_IWL<11550> A_IWL<11549> A_IWL<11548> A_IWL<11547> A_IWL<11546> A_IWL<11545> A_IWL<11544> A_IWL<11543> A_IWL<11542> A_IWL<11541> A_IWL<11540> A_IWL<11539> A_IWL<11538> A_IWL<11537> A_IWL<11536> A_IWL<11535> A_IWL<11534> A_IWL<11533> A_IWL<11532> A_IWL<11531> A_IWL<11530> A_IWL<11529> A_IWL<11528> A_IWL<11527> A_IWL<11526> A_IWL<11525> A_IWL<11524> A_IWL<11523> A_IWL<11522> A_IWL<11521> A_IWL<11520> A_IWL<11519> A_IWL<11518> A_IWL<11517> A_IWL<11516> A_IWL<11515> A_IWL<11514> A_IWL<11513> A_IWL<11512> A_IWL<11511> A_IWL<11510> A_IWL<11509> A_IWL<11508> A_IWL<11507> A_IWL<11506> A_IWL<11505> A_IWL<11504> A_IWL<11503> A_IWL<11502> A_IWL<11501> A_IWL<11500> A_IWL<11499> A_IWL<11498> A_IWL<11497> A_IWL<11496> A_IWL<11495> A_IWL<11494> A_IWL<11493> A_IWL<11492> A_IWL<11491> A_IWL<11490> A_IWL<11489> A_IWL<11488> A_IWL<11487> A_IWL<11486> A_IWL<11485> A_IWL<11484> A_IWL<11483> A_IWL<11482> A_IWL<11481> A_IWL<11480> A_IWL<11479> A_IWL<11478> A_IWL<11477> A_IWL<11476> A_IWL<11475> A_IWL<11474> A_IWL<11473> A_IWL<11472> A_IWL<11471> A_IWL<11470> A_IWL<11469> A_IWL<11468> A_IWL<11467> A_IWL<11466> A_IWL<11465> A_IWL<11464> A_IWL<11463> A_IWL<11462> A_IWL<11461> A_IWL<11460> A_IWL<11459> A_IWL<11458> A_IWL<11457> A_IWL<11456> A_IWL<11455> A_IWL<11454> A_IWL<11453> A_IWL<11452> A_IWL<11451> A_IWL<11450> A_IWL<11449> A_IWL<11448> A_IWL<11447> A_IWL<11446> A_IWL<11445> A_IWL<11444> A_IWL<11443> A_IWL<11442> A_IWL<11441> A_IWL<11440> A_IWL<11439> A_IWL<11438> A_IWL<11437> A_IWL<11436> A_IWL<11435> A_IWL<11434> A_IWL<11433> A_IWL<11432> A_IWL<11431> A_IWL<11430> A_IWL<11429> A_IWL<11428> A_IWL<11427> A_IWL<11426> A_IWL<11425> A_IWL<11424> A_IWL<11423> A_IWL<11422> A_IWL<11421> A_IWL<11420> A_IWL<11419> A_IWL<11418> A_IWL<11417> A_IWL<11416> A_IWL<11415> A_IWL<11414> A_IWL<11413> A_IWL<11412> A_IWL<11411> A_IWL<11410> A_IWL<11409> A_IWL<11408> A_IWL<11407> A_IWL<11406> A_IWL<11405> A_IWL<11404> A_IWL<11403> A_IWL<11402> A_IWL<11401> A_IWL<11400> A_IWL<11399> A_IWL<11398> A_IWL<11397> A_IWL<11396> A_IWL<11395> A_IWL<11394> A_IWL<11393> A_IWL<11392> A_IWL<11391> A_IWL<11390> A_IWL<11389> A_IWL<11388> A_IWL<11387> A_IWL<11386> A_IWL<11385> A_IWL<11384> A_IWL<11383> A_IWL<11382> A_IWL<11381> A_IWL<11380> A_IWL<11379> A_IWL<11378> A_IWL<11377> A_IWL<11376> A_IWL<11375> A_IWL<11374> A_IWL<11373> A_IWL<11372> A_IWL<11371> A_IWL<11370> A_IWL<11369> A_IWL<11368> A_IWL<11367> A_IWL<11366> A_IWL<11365> A_IWL<11364> A_IWL<11363> A_IWL<11362> A_IWL<11361> A_IWL<11360> A_IWL<11359> A_IWL<11358> A_IWL<11357> A_IWL<11356> A_IWL<11355> A_IWL<11354> A_IWL<11353> A_IWL<11352> A_IWL<11351> A_IWL<11350> A_IWL<11349> A_IWL<11348> A_IWL<11347> A_IWL<11346> A_IWL<11345> A_IWL<11344> A_IWL<11343> A_IWL<11342> A_IWL<11341> A_IWL<11340> A_IWL<11339> A_IWL<11338> A_IWL<11337> A_IWL<11336> A_IWL<11335> A_IWL<11334> A_IWL<11333> A_IWL<11332> A_IWL<11331> A_IWL<11330> A_IWL<11329> A_IWL<11328> A_IWL<11327> A_IWL<11326> A_IWL<11325> A_IWL<11324> A_IWL<11323> A_IWL<11322> A_IWL<11321> A_IWL<11320> A_IWL<11319> A_IWL<11318> A_IWL<11317> A_IWL<11316> A_IWL<11315> A_IWL<11314> A_IWL<11313> A_IWL<11312> A_IWL<11311> A_IWL<11310> A_IWL<11309> A_IWL<11308> A_IWL<11307> A_IWL<11306> A_IWL<11305> A_IWL<11304> A_IWL<11303> A_IWL<11302> A_IWL<11301> A_IWL<11300> A_IWL<11299> A_IWL<11298> A_IWL<11297> A_IWL<11296> A_IWL<11295> A_IWL<11294> A_IWL<11293> A_IWL<11292> A_IWL<11291> A_IWL<11290> A_IWL<11289> A_IWL<11288> A_IWL<11287> A_IWL<11286> A_IWL<11285> A_IWL<11284> A_IWL<11283> A_IWL<11282> A_IWL<11281> A_IWL<11280> A_IWL<11279> A_IWL<11278> A_IWL<11277> A_IWL<11276> A_IWL<11275> A_IWL<11274> A_IWL<11273> A_IWL<11272> A_IWL<11271> A_IWL<11270> A_IWL<11269> A_IWL<11268> A_IWL<11267> A_IWL<11266> A_IWL<11265> A_IWL<11264> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<21> A_BLC<43> A_BLC<42> A_BLC_TOP<43> A_BLC_TOP<42> A_BLT<43> A_BLT<42> A_BLT_TOP<43> A_BLT_TOP<42> A_IWL<10751> A_IWL<10750> A_IWL<10749> A_IWL<10748> A_IWL<10747> A_IWL<10746> A_IWL<10745> A_IWL<10744> A_IWL<10743> A_IWL<10742> A_IWL<10741> A_IWL<10740> A_IWL<10739> A_IWL<10738> A_IWL<10737> A_IWL<10736> A_IWL<10735> A_IWL<10734> A_IWL<10733> A_IWL<10732> A_IWL<10731> A_IWL<10730> A_IWL<10729> A_IWL<10728> A_IWL<10727> A_IWL<10726> A_IWL<10725> A_IWL<10724> A_IWL<10723> A_IWL<10722> A_IWL<10721> A_IWL<10720> A_IWL<10719> A_IWL<10718> A_IWL<10717> A_IWL<10716> A_IWL<10715> A_IWL<10714> A_IWL<10713> A_IWL<10712> A_IWL<10711> A_IWL<10710> A_IWL<10709> A_IWL<10708> A_IWL<10707> A_IWL<10706> A_IWL<10705> A_IWL<10704> A_IWL<10703> A_IWL<10702> A_IWL<10701> A_IWL<10700> A_IWL<10699> A_IWL<10698> A_IWL<10697> A_IWL<10696> A_IWL<10695> A_IWL<10694> A_IWL<10693> A_IWL<10692> A_IWL<10691> A_IWL<10690> A_IWL<10689> A_IWL<10688> A_IWL<10687> A_IWL<10686> A_IWL<10685> A_IWL<10684> A_IWL<10683> A_IWL<10682> A_IWL<10681> A_IWL<10680> A_IWL<10679> A_IWL<10678> A_IWL<10677> A_IWL<10676> A_IWL<10675> A_IWL<10674> A_IWL<10673> A_IWL<10672> A_IWL<10671> A_IWL<10670> A_IWL<10669> A_IWL<10668> A_IWL<10667> A_IWL<10666> A_IWL<10665> A_IWL<10664> A_IWL<10663> A_IWL<10662> A_IWL<10661> A_IWL<10660> A_IWL<10659> A_IWL<10658> A_IWL<10657> A_IWL<10656> A_IWL<10655> A_IWL<10654> A_IWL<10653> A_IWL<10652> A_IWL<10651> A_IWL<10650> A_IWL<10649> A_IWL<10648> A_IWL<10647> A_IWL<10646> A_IWL<10645> A_IWL<10644> A_IWL<10643> A_IWL<10642> A_IWL<10641> A_IWL<10640> A_IWL<10639> A_IWL<10638> A_IWL<10637> A_IWL<10636> A_IWL<10635> A_IWL<10634> A_IWL<10633> A_IWL<10632> A_IWL<10631> A_IWL<10630> A_IWL<10629> A_IWL<10628> A_IWL<10627> A_IWL<10626> A_IWL<10625> A_IWL<10624> A_IWL<10623> A_IWL<10622> A_IWL<10621> A_IWL<10620> A_IWL<10619> A_IWL<10618> A_IWL<10617> A_IWL<10616> A_IWL<10615> A_IWL<10614> A_IWL<10613> A_IWL<10612> A_IWL<10611> A_IWL<10610> A_IWL<10609> A_IWL<10608> A_IWL<10607> A_IWL<10606> A_IWL<10605> A_IWL<10604> A_IWL<10603> A_IWL<10602> A_IWL<10601> A_IWL<10600> A_IWL<10599> A_IWL<10598> A_IWL<10597> A_IWL<10596> A_IWL<10595> A_IWL<10594> A_IWL<10593> A_IWL<10592> A_IWL<10591> A_IWL<10590> A_IWL<10589> A_IWL<10588> A_IWL<10587> A_IWL<10586> A_IWL<10585> A_IWL<10584> A_IWL<10583> A_IWL<10582> A_IWL<10581> A_IWL<10580> A_IWL<10579> A_IWL<10578> A_IWL<10577> A_IWL<10576> A_IWL<10575> A_IWL<10574> A_IWL<10573> A_IWL<10572> A_IWL<10571> A_IWL<10570> A_IWL<10569> A_IWL<10568> A_IWL<10567> A_IWL<10566> A_IWL<10565> A_IWL<10564> A_IWL<10563> A_IWL<10562> A_IWL<10561> A_IWL<10560> A_IWL<10559> A_IWL<10558> A_IWL<10557> A_IWL<10556> A_IWL<10555> A_IWL<10554> A_IWL<10553> A_IWL<10552> A_IWL<10551> A_IWL<10550> A_IWL<10549> A_IWL<10548> A_IWL<10547> A_IWL<10546> A_IWL<10545> A_IWL<10544> A_IWL<10543> A_IWL<10542> A_IWL<10541> A_IWL<10540> A_IWL<10539> A_IWL<10538> A_IWL<10537> A_IWL<10536> A_IWL<10535> A_IWL<10534> A_IWL<10533> A_IWL<10532> A_IWL<10531> A_IWL<10530> A_IWL<10529> A_IWL<10528> A_IWL<10527> A_IWL<10526> A_IWL<10525> A_IWL<10524> A_IWL<10523> A_IWL<10522> A_IWL<10521> A_IWL<10520> A_IWL<10519> A_IWL<10518> A_IWL<10517> A_IWL<10516> A_IWL<10515> A_IWL<10514> A_IWL<10513> A_IWL<10512> A_IWL<10511> A_IWL<10510> A_IWL<10509> A_IWL<10508> A_IWL<10507> A_IWL<10506> A_IWL<10505> A_IWL<10504> A_IWL<10503> A_IWL<10502> A_IWL<10501> A_IWL<10500> A_IWL<10499> A_IWL<10498> A_IWL<10497> A_IWL<10496> A_IWL<10495> A_IWL<10494> A_IWL<10493> A_IWL<10492> A_IWL<10491> A_IWL<10490> A_IWL<10489> A_IWL<10488> A_IWL<10487> A_IWL<10486> A_IWL<10485> A_IWL<10484> A_IWL<10483> A_IWL<10482> A_IWL<10481> A_IWL<10480> A_IWL<10479> A_IWL<10478> A_IWL<10477> A_IWL<10476> A_IWL<10475> A_IWL<10474> A_IWL<10473> A_IWL<10472> A_IWL<10471> A_IWL<10470> A_IWL<10469> A_IWL<10468> A_IWL<10467> A_IWL<10466> A_IWL<10465> A_IWL<10464> A_IWL<10463> A_IWL<10462> A_IWL<10461> A_IWL<10460> A_IWL<10459> A_IWL<10458> A_IWL<10457> A_IWL<10456> A_IWL<10455> A_IWL<10454> A_IWL<10453> A_IWL<10452> A_IWL<10451> A_IWL<10450> A_IWL<10449> A_IWL<10448> A_IWL<10447> A_IWL<10446> A_IWL<10445> A_IWL<10444> A_IWL<10443> A_IWL<10442> A_IWL<10441> A_IWL<10440> A_IWL<10439> A_IWL<10438> A_IWL<10437> A_IWL<10436> A_IWL<10435> A_IWL<10434> A_IWL<10433> A_IWL<10432> A_IWL<10431> A_IWL<10430> A_IWL<10429> A_IWL<10428> A_IWL<10427> A_IWL<10426> A_IWL<10425> A_IWL<10424> A_IWL<10423> A_IWL<10422> A_IWL<10421> A_IWL<10420> A_IWL<10419> A_IWL<10418> A_IWL<10417> A_IWL<10416> A_IWL<10415> A_IWL<10414> A_IWL<10413> A_IWL<10412> A_IWL<10411> A_IWL<10410> A_IWL<10409> A_IWL<10408> A_IWL<10407> A_IWL<10406> A_IWL<10405> A_IWL<10404> A_IWL<10403> A_IWL<10402> A_IWL<10401> A_IWL<10400> A_IWL<10399> A_IWL<10398> A_IWL<10397> A_IWL<10396> A_IWL<10395> A_IWL<10394> A_IWL<10393> A_IWL<10392> A_IWL<10391> A_IWL<10390> A_IWL<10389> A_IWL<10388> A_IWL<10387> A_IWL<10386> A_IWL<10385> A_IWL<10384> A_IWL<10383> A_IWL<10382> A_IWL<10381> A_IWL<10380> A_IWL<10379> A_IWL<10378> A_IWL<10377> A_IWL<10376> A_IWL<10375> A_IWL<10374> A_IWL<10373> A_IWL<10372> A_IWL<10371> A_IWL<10370> A_IWL<10369> A_IWL<10368> A_IWL<10367> A_IWL<10366> A_IWL<10365> A_IWL<10364> A_IWL<10363> A_IWL<10362> A_IWL<10361> A_IWL<10360> A_IWL<10359> A_IWL<10358> A_IWL<10357> A_IWL<10356> A_IWL<10355> A_IWL<10354> A_IWL<10353> A_IWL<10352> A_IWL<10351> A_IWL<10350> A_IWL<10349> A_IWL<10348> A_IWL<10347> A_IWL<10346> A_IWL<10345> A_IWL<10344> A_IWL<10343> A_IWL<10342> A_IWL<10341> A_IWL<10340> A_IWL<10339> A_IWL<10338> A_IWL<10337> A_IWL<10336> A_IWL<10335> A_IWL<10334> A_IWL<10333> A_IWL<10332> A_IWL<10331> A_IWL<10330> A_IWL<10329> A_IWL<10328> A_IWL<10327> A_IWL<10326> A_IWL<10325> A_IWL<10324> A_IWL<10323> A_IWL<10322> A_IWL<10321> A_IWL<10320> A_IWL<10319> A_IWL<10318> A_IWL<10317> A_IWL<10316> A_IWL<10315> A_IWL<10314> A_IWL<10313> A_IWL<10312> A_IWL<10311> A_IWL<10310> A_IWL<10309> A_IWL<10308> A_IWL<10307> A_IWL<10306> A_IWL<10305> A_IWL<10304> A_IWL<10303> A_IWL<10302> A_IWL<10301> A_IWL<10300> A_IWL<10299> A_IWL<10298> A_IWL<10297> A_IWL<10296> A_IWL<10295> A_IWL<10294> A_IWL<10293> A_IWL<10292> A_IWL<10291> A_IWL<10290> A_IWL<10289> A_IWL<10288> A_IWL<10287> A_IWL<10286> A_IWL<10285> A_IWL<10284> A_IWL<10283> A_IWL<10282> A_IWL<10281> A_IWL<10280> A_IWL<10279> A_IWL<10278> A_IWL<10277> A_IWL<10276> A_IWL<10275> A_IWL<10274> A_IWL<10273> A_IWL<10272> A_IWL<10271> A_IWL<10270> A_IWL<10269> A_IWL<10268> A_IWL<10267> A_IWL<10266> A_IWL<10265> A_IWL<10264> A_IWL<10263> A_IWL<10262> A_IWL<10261> A_IWL<10260> A_IWL<10259> A_IWL<10258> A_IWL<10257> A_IWL<10256> A_IWL<10255> A_IWL<10254> A_IWL<10253> A_IWL<10252> A_IWL<10251> A_IWL<10250> A_IWL<10249> A_IWL<10248> A_IWL<10247> A_IWL<10246> A_IWL<10245> A_IWL<10244> A_IWL<10243> A_IWL<10242> A_IWL<10241> A_IWL<10240> A_IWL<11263> A_IWL<11262> A_IWL<11261> A_IWL<11260> A_IWL<11259> A_IWL<11258> A_IWL<11257> A_IWL<11256> A_IWL<11255> A_IWL<11254> A_IWL<11253> A_IWL<11252> A_IWL<11251> A_IWL<11250> A_IWL<11249> A_IWL<11248> A_IWL<11247> A_IWL<11246> A_IWL<11245> A_IWL<11244> A_IWL<11243> A_IWL<11242> A_IWL<11241> A_IWL<11240> A_IWL<11239> A_IWL<11238> A_IWL<11237> A_IWL<11236> A_IWL<11235> A_IWL<11234> A_IWL<11233> A_IWL<11232> A_IWL<11231> A_IWL<11230> A_IWL<11229> A_IWL<11228> A_IWL<11227> A_IWL<11226> A_IWL<11225> A_IWL<11224> A_IWL<11223> A_IWL<11222> A_IWL<11221> A_IWL<11220> A_IWL<11219> A_IWL<11218> A_IWL<11217> A_IWL<11216> A_IWL<11215> A_IWL<11214> A_IWL<11213> A_IWL<11212> A_IWL<11211> A_IWL<11210> A_IWL<11209> A_IWL<11208> A_IWL<11207> A_IWL<11206> A_IWL<11205> A_IWL<11204> A_IWL<11203> A_IWL<11202> A_IWL<11201> A_IWL<11200> A_IWL<11199> A_IWL<11198> A_IWL<11197> A_IWL<11196> A_IWL<11195> A_IWL<11194> A_IWL<11193> A_IWL<11192> A_IWL<11191> A_IWL<11190> A_IWL<11189> A_IWL<11188> A_IWL<11187> A_IWL<11186> A_IWL<11185> A_IWL<11184> A_IWL<11183> A_IWL<11182> A_IWL<11181> A_IWL<11180> A_IWL<11179> A_IWL<11178> A_IWL<11177> A_IWL<11176> A_IWL<11175> A_IWL<11174> A_IWL<11173> A_IWL<11172> A_IWL<11171> A_IWL<11170> A_IWL<11169> A_IWL<11168> A_IWL<11167> A_IWL<11166> A_IWL<11165> A_IWL<11164> A_IWL<11163> A_IWL<11162> A_IWL<11161> A_IWL<11160> A_IWL<11159> A_IWL<11158> A_IWL<11157> A_IWL<11156> A_IWL<11155> A_IWL<11154> A_IWL<11153> A_IWL<11152> A_IWL<11151> A_IWL<11150> A_IWL<11149> A_IWL<11148> A_IWL<11147> A_IWL<11146> A_IWL<11145> A_IWL<11144> A_IWL<11143> A_IWL<11142> A_IWL<11141> A_IWL<11140> A_IWL<11139> A_IWL<11138> A_IWL<11137> A_IWL<11136> A_IWL<11135> A_IWL<11134> A_IWL<11133> A_IWL<11132> A_IWL<11131> A_IWL<11130> A_IWL<11129> A_IWL<11128> A_IWL<11127> A_IWL<11126> A_IWL<11125> A_IWL<11124> A_IWL<11123> A_IWL<11122> A_IWL<11121> A_IWL<11120> A_IWL<11119> A_IWL<11118> A_IWL<11117> A_IWL<11116> A_IWL<11115> A_IWL<11114> A_IWL<11113> A_IWL<11112> A_IWL<11111> A_IWL<11110> A_IWL<11109> A_IWL<11108> A_IWL<11107> A_IWL<11106> A_IWL<11105> A_IWL<11104> A_IWL<11103> A_IWL<11102> A_IWL<11101> A_IWL<11100> A_IWL<11099> A_IWL<11098> A_IWL<11097> A_IWL<11096> A_IWL<11095> A_IWL<11094> A_IWL<11093> A_IWL<11092> A_IWL<11091> A_IWL<11090> A_IWL<11089> A_IWL<11088> A_IWL<11087> A_IWL<11086> A_IWL<11085> A_IWL<11084> A_IWL<11083> A_IWL<11082> A_IWL<11081> A_IWL<11080> A_IWL<11079> A_IWL<11078> A_IWL<11077> A_IWL<11076> A_IWL<11075> A_IWL<11074> A_IWL<11073> A_IWL<11072> A_IWL<11071> A_IWL<11070> A_IWL<11069> A_IWL<11068> A_IWL<11067> A_IWL<11066> A_IWL<11065> A_IWL<11064> A_IWL<11063> A_IWL<11062> A_IWL<11061> A_IWL<11060> A_IWL<11059> A_IWL<11058> A_IWL<11057> A_IWL<11056> A_IWL<11055> A_IWL<11054> A_IWL<11053> A_IWL<11052> A_IWL<11051> A_IWL<11050> A_IWL<11049> A_IWL<11048> A_IWL<11047> A_IWL<11046> A_IWL<11045> A_IWL<11044> A_IWL<11043> A_IWL<11042> A_IWL<11041> A_IWL<11040> A_IWL<11039> A_IWL<11038> A_IWL<11037> A_IWL<11036> A_IWL<11035> A_IWL<11034> A_IWL<11033> A_IWL<11032> A_IWL<11031> A_IWL<11030> A_IWL<11029> A_IWL<11028> A_IWL<11027> A_IWL<11026> A_IWL<11025> A_IWL<11024> A_IWL<11023> A_IWL<11022> A_IWL<11021> A_IWL<11020> A_IWL<11019> A_IWL<11018> A_IWL<11017> A_IWL<11016> A_IWL<11015> A_IWL<11014> A_IWL<11013> A_IWL<11012> A_IWL<11011> A_IWL<11010> A_IWL<11009> A_IWL<11008> A_IWL<11007> A_IWL<11006> A_IWL<11005> A_IWL<11004> A_IWL<11003> A_IWL<11002> A_IWL<11001> A_IWL<11000> A_IWL<10999> A_IWL<10998> A_IWL<10997> A_IWL<10996> A_IWL<10995> A_IWL<10994> A_IWL<10993> A_IWL<10992> A_IWL<10991> A_IWL<10990> A_IWL<10989> A_IWL<10988> A_IWL<10987> A_IWL<10986> A_IWL<10985> A_IWL<10984> A_IWL<10983> A_IWL<10982> A_IWL<10981> A_IWL<10980> A_IWL<10979> A_IWL<10978> A_IWL<10977> A_IWL<10976> A_IWL<10975> A_IWL<10974> A_IWL<10973> A_IWL<10972> A_IWL<10971> A_IWL<10970> A_IWL<10969> A_IWL<10968> A_IWL<10967> A_IWL<10966> A_IWL<10965> A_IWL<10964> A_IWL<10963> A_IWL<10962> A_IWL<10961> A_IWL<10960> A_IWL<10959> A_IWL<10958> A_IWL<10957> A_IWL<10956> A_IWL<10955> A_IWL<10954> A_IWL<10953> A_IWL<10952> A_IWL<10951> A_IWL<10950> A_IWL<10949> A_IWL<10948> A_IWL<10947> A_IWL<10946> A_IWL<10945> A_IWL<10944> A_IWL<10943> A_IWL<10942> A_IWL<10941> A_IWL<10940> A_IWL<10939> A_IWL<10938> A_IWL<10937> A_IWL<10936> A_IWL<10935> A_IWL<10934> A_IWL<10933> A_IWL<10932> A_IWL<10931> A_IWL<10930> A_IWL<10929> A_IWL<10928> A_IWL<10927> A_IWL<10926> A_IWL<10925> A_IWL<10924> A_IWL<10923> A_IWL<10922> A_IWL<10921> A_IWL<10920> A_IWL<10919> A_IWL<10918> A_IWL<10917> A_IWL<10916> A_IWL<10915> A_IWL<10914> A_IWL<10913> A_IWL<10912> A_IWL<10911> A_IWL<10910> A_IWL<10909> A_IWL<10908> A_IWL<10907> A_IWL<10906> A_IWL<10905> A_IWL<10904> A_IWL<10903> A_IWL<10902> A_IWL<10901> A_IWL<10900> A_IWL<10899> A_IWL<10898> A_IWL<10897> A_IWL<10896> A_IWL<10895> A_IWL<10894> A_IWL<10893> A_IWL<10892> A_IWL<10891> A_IWL<10890> A_IWL<10889> A_IWL<10888> A_IWL<10887> A_IWL<10886> A_IWL<10885> A_IWL<10884> A_IWL<10883> A_IWL<10882> A_IWL<10881> A_IWL<10880> A_IWL<10879> A_IWL<10878> A_IWL<10877> A_IWL<10876> A_IWL<10875> A_IWL<10874> A_IWL<10873> A_IWL<10872> A_IWL<10871> A_IWL<10870> A_IWL<10869> A_IWL<10868> A_IWL<10867> A_IWL<10866> A_IWL<10865> A_IWL<10864> A_IWL<10863> A_IWL<10862> A_IWL<10861> A_IWL<10860> A_IWL<10859> A_IWL<10858> A_IWL<10857> A_IWL<10856> A_IWL<10855> A_IWL<10854> A_IWL<10853> A_IWL<10852> A_IWL<10851> A_IWL<10850> A_IWL<10849> A_IWL<10848> A_IWL<10847> A_IWL<10846> A_IWL<10845> A_IWL<10844> A_IWL<10843> A_IWL<10842> A_IWL<10841> A_IWL<10840> A_IWL<10839> A_IWL<10838> A_IWL<10837> A_IWL<10836> A_IWL<10835> A_IWL<10834> A_IWL<10833> A_IWL<10832> A_IWL<10831> A_IWL<10830> A_IWL<10829> A_IWL<10828> A_IWL<10827> A_IWL<10826> A_IWL<10825> A_IWL<10824> A_IWL<10823> A_IWL<10822> A_IWL<10821> A_IWL<10820> A_IWL<10819> A_IWL<10818> A_IWL<10817> A_IWL<10816> A_IWL<10815> A_IWL<10814> A_IWL<10813> A_IWL<10812> A_IWL<10811> A_IWL<10810> A_IWL<10809> A_IWL<10808> A_IWL<10807> A_IWL<10806> A_IWL<10805> A_IWL<10804> A_IWL<10803> A_IWL<10802> A_IWL<10801> A_IWL<10800> A_IWL<10799> A_IWL<10798> A_IWL<10797> A_IWL<10796> A_IWL<10795> A_IWL<10794> A_IWL<10793> A_IWL<10792> A_IWL<10791> A_IWL<10790> A_IWL<10789> A_IWL<10788> A_IWL<10787> A_IWL<10786> A_IWL<10785> A_IWL<10784> A_IWL<10783> A_IWL<10782> A_IWL<10781> A_IWL<10780> A_IWL<10779> A_IWL<10778> A_IWL<10777> A_IWL<10776> A_IWL<10775> A_IWL<10774> A_IWL<10773> A_IWL<10772> A_IWL<10771> A_IWL<10770> A_IWL<10769> A_IWL<10768> A_IWL<10767> A_IWL<10766> A_IWL<10765> A_IWL<10764> A_IWL<10763> A_IWL<10762> A_IWL<10761> A_IWL<10760> A_IWL<10759> A_IWL<10758> A_IWL<10757> A_IWL<10756> A_IWL<10755> A_IWL<10754> A_IWL<10753> A_IWL<10752> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<20> A_BLC<41> A_BLC<40> A_BLC_TOP<41> A_BLC_TOP<40> A_BLT<41> A_BLT<40> A_BLT_TOP<41> A_BLT_TOP<40> A_IWL<10239> A_IWL<10238> A_IWL<10237> A_IWL<10236> A_IWL<10235> A_IWL<10234> A_IWL<10233> A_IWL<10232> A_IWL<10231> A_IWL<10230> A_IWL<10229> A_IWL<10228> A_IWL<10227> A_IWL<10226> A_IWL<10225> A_IWL<10224> A_IWL<10223> A_IWL<10222> A_IWL<10221> A_IWL<10220> A_IWL<10219> A_IWL<10218> A_IWL<10217> A_IWL<10216> A_IWL<10215> A_IWL<10214> A_IWL<10213> A_IWL<10212> A_IWL<10211> A_IWL<10210> A_IWL<10209> A_IWL<10208> A_IWL<10207> A_IWL<10206> A_IWL<10205> A_IWL<10204> A_IWL<10203> A_IWL<10202> A_IWL<10201> A_IWL<10200> A_IWL<10199> A_IWL<10198> A_IWL<10197> A_IWL<10196> A_IWL<10195> A_IWL<10194> A_IWL<10193> A_IWL<10192> A_IWL<10191> A_IWL<10190> A_IWL<10189> A_IWL<10188> A_IWL<10187> A_IWL<10186> A_IWL<10185> A_IWL<10184> A_IWL<10183> A_IWL<10182> A_IWL<10181> A_IWL<10180> A_IWL<10179> A_IWL<10178> A_IWL<10177> A_IWL<10176> A_IWL<10175> A_IWL<10174> A_IWL<10173> A_IWL<10172> A_IWL<10171> A_IWL<10170> A_IWL<10169> A_IWL<10168> A_IWL<10167> A_IWL<10166> A_IWL<10165> A_IWL<10164> A_IWL<10163> A_IWL<10162> A_IWL<10161> A_IWL<10160> A_IWL<10159> A_IWL<10158> A_IWL<10157> A_IWL<10156> A_IWL<10155> A_IWL<10154> A_IWL<10153> A_IWL<10152> A_IWL<10151> A_IWL<10150> A_IWL<10149> A_IWL<10148> A_IWL<10147> A_IWL<10146> A_IWL<10145> A_IWL<10144> A_IWL<10143> A_IWL<10142> A_IWL<10141> A_IWL<10140> A_IWL<10139> A_IWL<10138> A_IWL<10137> A_IWL<10136> A_IWL<10135> A_IWL<10134> A_IWL<10133> A_IWL<10132> A_IWL<10131> A_IWL<10130> A_IWL<10129> A_IWL<10128> A_IWL<10127> A_IWL<10126> A_IWL<10125> A_IWL<10124> A_IWL<10123> A_IWL<10122> A_IWL<10121> A_IWL<10120> A_IWL<10119> A_IWL<10118> A_IWL<10117> A_IWL<10116> A_IWL<10115> A_IWL<10114> A_IWL<10113> A_IWL<10112> A_IWL<10111> A_IWL<10110> A_IWL<10109> A_IWL<10108> A_IWL<10107> A_IWL<10106> A_IWL<10105> A_IWL<10104> A_IWL<10103> A_IWL<10102> A_IWL<10101> A_IWL<10100> A_IWL<10099> A_IWL<10098> A_IWL<10097> A_IWL<10096> A_IWL<10095> A_IWL<10094> A_IWL<10093> A_IWL<10092> A_IWL<10091> A_IWL<10090> A_IWL<10089> A_IWL<10088> A_IWL<10087> A_IWL<10086> A_IWL<10085> A_IWL<10084> A_IWL<10083> A_IWL<10082> A_IWL<10081> A_IWL<10080> A_IWL<10079> A_IWL<10078> A_IWL<10077> A_IWL<10076> A_IWL<10075> A_IWL<10074> A_IWL<10073> A_IWL<10072> A_IWL<10071> A_IWL<10070> A_IWL<10069> A_IWL<10068> A_IWL<10067> A_IWL<10066> A_IWL<10065> A_IWL<10064> A_IWL<10063> A_IWL<10062> A_IWL<10061> A_IWL<10060> A_IWL<10059> A_IWL<10058> A_IWL<10057> A_IWL<10056> A_IWL<10055> A_IWL<10054> A_IWL<10053> A_IWL<10052> A_IWL<10051> A_IWL<10050> A_IWL<10049> A_IWL<10048> A_IWL<10047> A_IWL<10046> A_IWL<10045> A_IWL<10044> A_IWL<10043> A_IWL<10042> A_IWL<10041> A_IWL<10040> A_IWL<10039> A_IWL<10038> A_IWL<10037> A_IWL<10036> A_IWL<10035> A_IWL<10034> A_IWL<10033> A_IWL<10032> A_IWL<10031> A_IWL<10030> A_IWL<10029> A_IWL<10028> A_IWL<10027> A_IWL<10026> A_IWL<10025> A_IWL<10024> A_IWL<10023> A_IWL<10022> A_IWL<10021> A_IWL<10020> A_IWL<10019> A_IWL<10018> A_IWL<10017> A_IWL<10016> A_IWL<10015> A_IWL<10014> A_IWL<10013> A_IWL<10012> A_IWL<10011> A_IWL<10010> A_IWL<10009> A_IWL<10008> A_IWL<10007> A_IWL<10006> A_IWL<10005> A_IWL<10004> A_IWL<10003> A_IWL<10002> A_IWL<10001> A_IWL<10000> A_IWL<9999> A_IWL<9998> A_IWL<9997> A_IWL<9996> A_IWL<9995> A_IWL<9994> A_IWL<9993> A_IWL<9992> A_IWL<9991> A_IWL<9990> A_IWL<9989> A_IWL<9988> A_IWL<9987> A_IWL<9986> A_IWL<9985> A_IWL<9984> A_IWL<9983> A_IWL<9982> A_IWL<9981> A_IWL<9980> A_IWL<9979> A_IWL<9978> A_IWL<9977> A_IWL<9976> A_IWL<9975> A_IWL<9974> A_IWL<9973> A_IWL<9972> A_IWL<9971> A_IWL<9970> A_IWL<9969> A_IWL<9968> A_IWL<9967> A_IWL<9966> A_IWL<9965> A_IWL<9964> A_IWL<9963> A_IWL<9962> A_IWL<9961> A_IWL<9960> A_IWL<9959> A_IWL<9958> A_IWL<9957> A_IWL<9956> A_IWL<9955> A_IWL<9954> A_IWL<9953> A_IWL<9952> A_IWL<9951> A_IWL<9950> A_IWL<9949> A_IWL<9948> A_IWL<9947> A_IWL<9946> A_IWL<9945> A_IWL<9944> A_IWL<9943> A_IWL<9942> A_IWL<9941> A_IWL<9940> A_IWL<9939> A_IWL<9938> A_IWL<9937> A_IWL<9936> A_IWL<9935> A_IWL<9934> A_IWL<9933> A_IWL<9932> A_IWL<9931> A_IWL<9930> A_IWL<9929> A_IWL<9928> A_IWL<9927> A_IWL<9926> A_IWL<9925> A_IWL<9924> A_IWL<9923> A_IWL<9922> A_IWL<9921> A_IWL<9920> A_IWL<9919> A_IWL<9918> A_IWL<9917> A_IWL<9916> A_IWL<9915> A_IWL<9914> A_IWL<9913> A_IWL<9912> A_IWL<9911> A_IWL<9910> A_IWL<9909> A_IWL<9908> A_IWL<9907> A_IWL<9906> A_IWL<9905> A_IWL<9904> A_IWL<9903> A_IWL<9902> A_IWL<9901> A_IWL<9900> A_IWL<9899> A_IWL<9898> A_IWL<9897> A_IWL<9896> A_IWL<9895> A_IWL<9894> A_IWL<9893> A_IWL<9892> A_IWL<9891> A_IWL<9890> A_IWL<9889> A_IWL<9888> A_IWL<9887> A_IWL<9886> A_IWL<9885> A_IWL<9884> A_IWL<9883> A_IWL<9882> A_IWL<9881> A_IWL<9880> A_IWL<9879> A_IWL<9878> A_IWL<9877> A_IWL<9876> A_IWL<9875> A_IWL<9874> A_IWL<9873> A_IWL<9872> A_IWL<9871> A_IWL<9870> A_IWL<9869> A_IWL<9868> A_IWL<9867> A_IWL<9866> A_IWL<9865> A_IWL<9864> A_IWL<9863> A_IWL<9862> A_IWL<9861> A_IWL<9860> A_IWL<9859> A_IWL<9858> A_IWL<9857> A_IWL<9856> A_IWL<9855> A_IWL<9854> A_IWL<9853> A_IWL<9852> A_IWL<9851> A_IWL<9850> A_IWL<9849> A_IWL<9848> A_IWL<9847> A_IWL<9846> A_IWL<9845> A_IWL<9844> A_IWL<9843> A_IWL<9842> A_IWL<9841> A_IWL<9840> A_IWL<9839> A_IWL<9838> A_IWL<9837> A_IWL<9836> A_IWL<9835> A_IWL<9834> A_IWL<9833> A_IWL<9832> A_IWL<9831> A_IWL<9830> A_IWL<9829> A_IWL<9828> A_IWL<9827> A_IWL<9826> A_IWL<9825> A_IWL<9824> A_IWL<9823> A_IWL<9822> A_IWL<9821> A_IWL<9820> A_IWL<9819> A_IWL<9818> A_IWL<9817> A_IWL<9816> A_IWL<9815> A_IWL<9814> A_IWL<9813> A_IWL<9812> A_IWL<9811> A_IWL<9810> A_IWL<9809> A_IWL<9808> A_IWL<9807> A_IWL<9806> A_IWL<9805> A_IWL<9804> A_IWL<9803> A_IWL<9802> A_IWL<9801> A_IWL<9800> A_IWL<9799> A_IWL<9798> A_IWL<9797> A_IWL<9796> A_IWL<9795> A_IWL<9794> A_IWL<9793> A_IWL<9792> A_IWL<9791> A_IWL<9790> A_IWL<9789> A_IWL<9788> A_IWL<9787> A_IWL<9786> A_IWL<9785> A_IWL<9784> A_IWL<9783> A_IWL<9782> A_IWL<9781> A_IWL<9780> A_IWL<9779> A_IWL<9778> A_IWL<9777> A_IWL<9776> A_IWL<9775> A_IWL<9774> A_IWL<9773> A_IWL<9772> A_IWL<9771> A_IWL<9770> A_IWL<9769> A_IWL<9768> A_IWL<9767> A_IWL<9766> A_IWL<9765> A_IWL<9764> A_IWL<9763> A_IWL<9762> A_IWL<9761> A_IWL<9760> A_IWL<9759> A_IWL<9758> A_IWL<9757> A_IWL<9756> A_IWL<9755> A_IWL<9754> A_IWL<9753> A_IWL<9752> A_IWL<9751> A_IWL<9750> A_IWL<9749> A_IWL<9748> A_IWL<9747> A_IWL<9746> A_IWL<9745> A_IWL<9744> A_IWL<9743> A_IWL<9742> A_IWL<9741> A_IWL<9740> A_IWL<9739> A_IWL<9738> A_IWL<9737> A_IWL<9736> A_IWL<9735> A_IWL<9734> A_IWL<9733> A_IWL<9732> A_IWL<9731> A_IWL<9730> A_IWL<9729> A_IWL<9728> A_IWL<10751> A_IWL<10750> A_IWL<10749> A_IWL<10748> A_IWL<10747> A_IWL<10746> A_IWL<10745> A_IWL<10744> A_IWL<10743> A_IWL<10742> A_IWL<10741> A_IWL<10740> A_IWL<10739> A_IWL<10738> A_IWL<10737> A_IWL<10736> A_IWL<10735> A_IWL<10734> A_IWL<10733> A_IWL<10732> A_IWL<10731> A_IWL<10730> A_IWL<10729> A_IWL<10728> A_IWL<10727> A_IWL<10726> A_IWL<10725> A_IWL<10724> A_IWL<10723> A_IWL<10722> A_IWL<10721> A_IWL<10720> A_IWL<10719> A_IWL<10718> A_IWL<10717> A_IWL<10716> A_IWL<10715> A_IWL<10714> A_IWL<10713> A_IWL<10712> A_IWL<10711> A_IWL<10710> A_IWL<10709> A_IWL<10708> A_IWL<10707> A_IWL<10706> A_IWL<10705> A_IWL<10704> A_IWL<10703> A_IWL<10702> A_IWL<10701> A_IWL<10700> A_IWL<10699> A_IWL<10698> A_IWL<10697> A_IWL<10696> A_IWL<10695> A_IWL<10694> A_IWL<10693> A_IWL<10692> A_IWL<10691> A_IWL<10690> A_IWL<10689> A_IWL<10688> A_IWL<10687> A_IWL<10686> A_IWL<10685> A_IWL<10684> A_IWL<10683> A_IWL<10682> A_IWL<10681> A_IWL<10680> A_IWL<10679> A_IWL<10678> A_IWL<10677> A_IWL<10676> A_IWL<10675> A_IWL<10674> A_IWL<10673> A_IWL<10672> A_IWL<10671> A_IWL<10670> A_IWL<10669> A_IWL<10668> A_IWL<10667> A_IWL<10666> A_IWL<10665> A_IWL<10664> A_IWL<10663> A_IWL<10662> A_IWL<10661> A_IWL<10660> A_IWL<10659> A_IWL<10658> A_IWL<10657> A_IWL<10656> A_IWL<10655> A_IWL<10654> A_IWL<10653> A_IWL<10652> A_IWL<10651> A_IWL<10650> A_IWL<10649> A_IWL<10648> A_IWL<10647> A_IWL<10646> A_IWL<10645> A_IWL<10644> A_IWL<10643> A_IWL<10642> A_IWL<10641> A_IWL<10640> A_IWL<10639> A_IWL<10638> A_IWL<10637> A_IWL<10636> A_IWL<10635> A_IWL<10634> A_IWL<10633> A_IWL<10632> A_IWL<10631> A_IWL<10630> A_IWL<10629> A_IWL<10628> A_IWL<10627> A_IWL<10626> A_IWL<10625> A_IWL<10624> A_IWL<10623> A_IWL<10622> A_IWL<10621> A_IWL<10620> A_IWL<10619> A_IWL<10618> A_IWL<10617> A_IWL<10616> A_IWL<10615> A_IWL<10614> A_IWL<10613> A_IWL<10612> A_IWL<10611> A_IWL<10610> A_IWL<10609> A_IWL<10608> A_IWL<10607> A_IWL<10606> A_IWL<10605> A_IWL<10604> A_IWL<10603> A_IWL<10602> A_IWL<10601> A_IWL<10600> A_IWL<10599> A_IWL<10598> A_IWL<10597> A_IWL<10596> A_IWL<10595> A_IWL<10594> A_IWL<10593> A_IWL<10592> A_IWL<10591> A_IWL<10590> A_IWL<10589> A_IWL<10588> A_IWL<10587> A_IWL<10586> A_IWL<10585> A_IWL<10584> A_IWL<10583> A_IWL<10582> A_IWL<10581> A_IWL<10580> A_IWL<10579> A_IWL<10578> A_IWL<10577> A_IWL<10576> A_IWL<10575> A_IWL<10574> A_IWL<10573> A_IWL<10572> A_IWL<10571> A_IWL<10570> A_IWL<10569> A_IWL<10568> A_IWL<10567> A_IWL<10566> A_IWL<10565> A_IWL<10564> A_IWL<10563> A_IWL<10562> A_IWL<10561> A_IWL<10560> A_IWL<10559> A_IWL<10558> A_IWL<10557> A_IWL<10556> A_IWL<10555> A_IWL<10554> A_IWL<10553> A_IWL<10552> A_IWL<10551> A_IWL<10550> A_IWL<10549> A_IWL<10548> A_IWL<10547> A_IWL<10546> A_IWL<10545> A_IWL<10544> A_IWL<10543> A_IWL<10542> A_IWL<10541> A_IWL<10540> A_IWL<10539> A_IWL<10538> A_IWL<10537> A_IWL<10536> A_IWL<10535> A_IWL<10534> A_IWL<10533> A_IWL<10532> A_IWL<10531> A_IWL<10530> A_IWL<10529> A_IWL<10528> A_IWL<10527> A_IWL<10526> A_IWL<10525> A_IWL<10524> A_IWL<10523> A_IWL<10522> A_IWL<10521> A_IWL<10520> A_IWL<10519> A_IWL<10518> A_IWL<10517> A_IWL<10516> A_IWL<10515> A_IWL<10514> A_IWL<10513> A_IWL<10512> A_IWL<10511> A_IWL<10510> A_IWL<10509> A_IWL<10508> A_IWL<10507> A_IWL<10506> A_IWL<10505> A_IWL<10504> A_IWL<10503> A_IWL<10502> A_IWL<10501> A_IWL<10500> A_IWL<10499> A_IWL<10498> A_IWL<10497> A_IWL<10496> A_IWL<10495> A_IWL<10494> A_IWL<10493> A_IWL<10492> A_IWL<10491> A_IWL<10490> A_IWL<10489> A_IWL<10488> A_IWL<10487> A_IWL<10486> A_IWL<10485> A_IWL<10484> A_IWL<10483> A_IWL<10482> A_IWL<10481> A_IWL<10480> A_IWL<10479> A_IWL<10478> A_IWL<10477> A_IWL<10476> A_IWL<10475> A_IWL<10474> A_IWL<10473> A_IWL<10472> A_IWL<10471> A_IWL<10470> A_IWL<10469> A_IWL<10468> A_IWL<10467> A_IWL<10466> A_IWL<10465> A_IWL<10464> A_IWL<10463> A_IWL<10462> A_IWL<10461> A_IWL<10460> A_IWL<10459> A_IWL<10458> A_IWL<10457> A_IWL<10456> A_IWL<10455> A_IWL<10454> A_IWL<10453> A_IWL<10452> A_IWL<10451> A_IWL<10450> A_IWL<10449> A_IWL<10448> A_IWL<10447> A_IWL<10446> A_IWL<10445> A_IWL<10444> A_IWL<10443> A_IWL<10442> A_IWL<10441> A_IWL<10440> A_IWL<10439> A_IWL<10438> A_IWL<10437> A_IWL<10436> A_IWL<10435> A_IWL<10434> A_IWL<10433> A_IWL<10432> A_IWL<10431> A_IWL<10430> A_IWL<10429> A_IWL<10428> A_IWL<10427> A_IWL<10426> A_IWL<10425> A_IWL<10424> A_IWL<10423> A_IWL<10422> A_IWL<10421> A_IWL<10420> A_IWL<10419> A_IWL<10418> A_IWL<10417> A_IWL<10416> A_IWL<10415> A_IWL<10414> A_IWL<10413> A_IWL<10412> A_IWL<10411> A_IWL<10410> A_IWL<10409> A_IWL<10408> A_IWL<10407> A_IWL<10406> A_IWL<10405> A_IWL<10404> A_IWL<10403> A_IWL<10402> A_IWL<10401> A_IWL<10400> A_IWL<10399> A_IWL<10398> A_IWL<10397> A_IWL<10396> A_IWL<10395> A_IWL<10394> A_IWL<10393> A_IWL<10392> A_IWL<10391> A_IWL<10390> A_IWL<10389> A_IWL<10388> A_IWL<10387> A_IWL<10386> A_IWL<10385> A_IWL<10384> A_IWL<10383> A_IWL<10382> A_IWL<10381> A_IWL<10380> A_IWL<10379> A_IWL<10378> A_IWL<10377> A_IWL<10376> A_IWL<10375> A_IWL<10374> A_IWL<10373> A_IWL<10372> A_IWL<10371> A_IWL<10370> A_IWL<10369> A_IWL<10368> A_IWL<10367> A_IWL<10366> A_IWL<10365> A_IWL<10364> A_IWL<10363> A_IWL<10362> A_IWL<10361> A_IWL<10360> A_IWL<10359> A_IWL<10358> A_IWL<10357> A_IWL<10356> A_IWL<10355> A_IWL<10354> A_IWL<10353> A_IWL<10352> A_IWL<10351> A_IWL<10350> A_IWL<10349> A_IWL<10348> A_IWL<10347> A_IWL<10346> A_IWL<10345> A_IWL<10344> A_IWL<10343> A_IWL<10342> A_IWL<10341> A_IWL<10340> A_IWL<10339> A_IWL<10338> A_IWL<10337> A_IWL<10336> A_IWL<10335> A_IWL<10334> A_IWL<10333> A_IWL<10332> A_IWL<10331> A_IWL<10330> A_IWL<10329> A_IWL<10328> A_IWL<10327> A_IWL<10326> A_IWL<10325> A_IWL<10324> A_IWL<10323> A_IWL<10322> A_IWL<10321> A_IWL<10320> A_IWL<10319> A_IWL<10318> A_IWL<10317> A_IWL<10316> A_IWL<10315> A_IWL<10314> A_IWL<10313> A_IWL<10312> A_IWL<10311> A_IWL<10310> A_IWL<10309> A_IWL<10308> A_IWL<10307> A_IWL<10306> A_IWL<10305> A_IWL<10304> A_IWL<10303> A_IWL<10302> A_IWL<10301> A_IWL<10300> A_IWL<10299> A_IWL<10298> A_IWL<10297> A_IWL<10296> A_IWL<10295> A_IWL<10294> A_IWL<10293> A_IWL<10292> A_IWL<10291> A_IWL<10290> A_IWL<10289> A_IWL<10288> A_IWL<10287> A_IWL<10286> A_IWL<10285> A_IWL<10284> A_IWL<10283> A_IWL<10282> A_IWL<10281> A_IWL<10280> A_IWL<10279> A_IWL<10278> A_IWL<10277> A_IWL<10276> A_IWL<10275> A_IWL<10274> A_IWL<10273> A_IWL<10272> A_IWL<10271> A_IWL<10270> A_IWL<10269> A_IWL<10268> A_IWL<10267> A_IWL<10266> A_IWL<10265> A_IWL<10264> A_IWL<10263> A_IWL<10262> A_IWL<10261> A_IWL<10260> A_IWL<10259> A_IWL<10258> A_IWL<10257> A_IWL<10256> A_IWL<10255> A_IWL<10254> A_IWL<10253> A_IWL<10252> A_IWL<10251> A_IWL<10250> A_IWL<10249> A_IWL<10248> A_IWL<10247> A_IWL<10246> A_IWL<10245> A_IWL<10244> A_IWL<10243> A_IWL<10242> A_IWL<10241> A_IWL<10240> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<19> A_BLC<39> A_BLC<38> A_BLC_TOP<39> A_BLC_TOP<38> A_BLT<39> A_BLT<38> A_BLT_TOP<39> A_BLT_TOP<38> A_IWL<9727> A_IWL<9726> A_IWL<9725> A_IWL<9724> A_IWL<9723> A_IWL<9722> A_IWL<9721> A_IWL<9720> A_IWL<9719> A_IWL<9718> A_IWL<9717> A_IWL<9716> A_IWL<9715> A_IWL<9714> A_IWL<9713> A_IWL<9712> A_IWL<9711> A_IWL<9710> A_IWL<9709> A_IWL<9708> A_IWL<9707> A_IWL<9706> A_IWL<9705> A_IWL<9704> A_IWL<9703> A_IWL<9702> A_IWL<9701> A_IWL<9700> A_IWL<9699> A_IWL<9698> A_IWL<9697> A_IWL<9696> A_IWL<9695> A_IWL<9694> A_IWL<9693> A_IWL<9692> A_IWL<9691> A_IWL<9690> A_IWL<9689> A_IWL<9688> A_IWL<9687> A_IWL<9686> A_IWL<9685> A_IWL<9684> A_IWL<9683> A_IWL<9682> A_IWL<9681> A_IWL<9680> A_IWL<9679> A_IWL<9678> A_IWL<9677> A_IWL<9676> A_IWL<9675> A_IWL<9674> A_IWL<9673> A_IWL<9672> A_IWL<9671> A_IWL<9670> A_IWL<9669> A_IWL<9668> A_IWL<9667> A_IWL<9666> A_IWL<9665> A_IWL<9664> A_IWL<9663> A_IWL<9662> A_IWL<9661> A_IWL<9660> A_IWL<9659> A_IWL<9658> A_IWL<9657> A_IWL<9656> A_IWL<9655> A_IWL<9654> A_IWL<9653> A_IWL<9652> A_IWL<9651> A_IWL<9650> A_IWL<9649> A_IWL<9648> A_IWL<9647> A_IWL<9646> A_IWL<9645> A_IWL<9644> A_IWL<9643> A_IWL<9642> A_IWL<9641> A_IWL<9640> A_IWL<9639> A_IWL<9638> A_IWL<9637> A_IWL<9636> A_IWL<9635> A_IWL<9634> A_IWL<9633> A_IWL<9632> A_IWL<9631> A_IWL<9630> A_IWL<9629> A_IWL<9628> A_IWL<9627> A_IWL<9626> A_IWL<9625> A_IWL<9624> A_IWL<9623> A_IWL<9622> A_IWL<9621> A_IWL<9620> A_IWL<9619> A_IWL<9618> A_IWL<9617> A_IWL<9616> A_IWL<9615> A_IWL<9614> A_IWL<9613> A_IWL<9612> A_IWL<9611> A_IWL<9610> A_IWL<9609> A_IWL<9608> A_IWL<9607> A_IWL<9606> A_IWL<9605> A_IWL<9604> A_IWL<9603> A_IWL<9602> A_IWL<9601> A_IWL<9600> A_IWL<9599> A_IWL<9598> A_IWL<9597> A_IWL<9596> A_IWL<9595> A_IWL<9594> A_IWL<9593> A_IWL<9592> A_IWL<9591> A_IWL<9590> A_IWL<9589> A_IWL<9588> A_IWL<9587> A_IWL<9586> A_IWL<9585> A_IWL<9584> A_IWL<9583> A_IWL<9582> A_IWL<9581> A_IWL<9580> A_IWL<9579> A_IWL<9578> A_IWL<9577> A_IWL<9576> A_IWL<9575> A_IWL<9574> A_IWL<9573> A_IWL<9572> A_IWL<9571> A_IWL<9570> A_IWL<9569> A_IWL<9568> A_IWL<9567> A_IWL<9566> A_IWL<9565> A_IWL<9564> A_IWL<9563> A_IWL<9562> A_IWL<9561> A_IWL<9560> A_IWL<9559> A_IWL<9558> A_IWL<9557> A_IWL<9556> A_IWL<9555> A_IWL<9554> A_IWL<9553> A_IWL<9552> A_IWL<9551> A_IWL<9550> A_IWL<9549> A_IWL<9548> A_IWL<9547> A_IWL<9546> A_IWL<9545> A_IWL<9544> A_IWL<9543> A_IWL<9542> A_IWL<9541> A_IWL<9540> A_IWL<9539> A_IWL<9538> A_IWL<9537> A_IWL<9536> A_IWL<9535> A_IWL<9534> A_IWL<9533> A_IWL<9532> A_IWL<9531> A_IWL<9530> A_IWL<9529> A_IWL<9528> A_IWL<9527> A_IWL<9526> A_IWL<9525> A_IWL<9524> A_IWL<9523> A_IWL<9522> A_IWL<9521> A_IWL<9520> A_IWL<9519> A_IWL<9518> A_IWL<9517> A_IWL<9516> A_IWL<9515> A_IWL<9514> A_IWL<9513> A_IWL<9512> A_IWL<9511> A_IWL<9510> A_IWL<9509> A_IWL<9508> A_IWL<9507> A_IWL<9506> A_IWL<9505> A_IWL<9504> A_IWL<9503> A_IWL<9502> A_IWL<9501> A_IWL<9500> A_IWL<9499> A_IWL<9498> A_IWL<9497> A_IWL<9496> A_IWL<9495> A_IWL<9494> A_IWL<9493> A_IWL<9492> A_IWL<9491> A_IWL<9490> A_IWL<9489> A_IWL<9488> A_IWL<9487> A_IWL<9486> A_IWL<9485> A_IWL<9484> A_IWL<9483> A_IWL<9482> A_IWL<9481> A_IWL<9480> A_IWL<9479> A_IWL<9478> A_IWL<9477> A_IWL<9476> A_IWL<9475> A_IWL<9474> A_IWL<9473> A_IWL<9472> A_IWL<9471> A_IWL<9470> A_IWL<9469> A_IWL<9468> A_IWL<9467> A_IWL<9466> A_IWL<9465> A_IWL<9464> A_IWL<9463> A_IWL<9462> A_IWL<9461> A_IWL<9460> A_IWL<9459> A_IWL<9458> A_IWL<9457> A_IWL<9456> A_IWL<9455> A_IWL<9454> A_IWL<9453> A_IWL<9452> A_IWL<9451> A_IWL<9450> A_IWL<9449> A_IWL<9448> A_IWL<9447> A_IWL<9446> A_IWL<9445> A_IWL<9444> A_IWL<9443> A_IWL<9442> A_IWL<9441> A_IWL<9440> A_IWL<9439> A_IWL<9438> A_IWL<9437> A_IWL<9436> A_IWL<9435> A_IWL<9434> A_IWL<9433> A_IWL<9432> A_IWL<9431> A_IWL<9430> A_IWL<9429> A_IWL<9428> A_IWL<9427> A_IWL<9426> A_IWL<9425> A_IWL<9424> A_IWL<9423> A_IWL<9422> A_IWL<9421> A_IWL<9420> A_IWL<9419> A_IWL<9418> A_IWL<9417> A_IWL<9416> A_IWL<9415> A_IWL<9414> A_IWL<9413> A_IWL<9412> A_IWL<9411> A_IWL<9410> A_IWL<9409> A_IWL<9408> A_IWL<9407> A_IWL<9406> A_IWL<9405> A_IWL<9404> A_IWL<9403> A_IWL<9402> A_IWL<9401> A_IWL<9400> A_IWL<9399> A_IWL<9398> A_IWL<9397> A_IWL<9396> A_IWL<9395> A_IWL<9394> A_IWL<9393> A_IWL<9392> A_IWL<9391> A_IWL<9390> A_IWL<9389> A_IWL<9388> A_IWL<9387> A_IWL<9386> A_IWL<9385> A_IWL<9384> A_IWL<9383> A_IWL<9382> A_IWL<9381> A_IWL<9380> A_IWL<9379> A_IWL<9378> A_IWL<9377> A_IWL<9376> A_IWL<9375> A_IWL<9374> A_IWL<9373> A_IWL<9372> A_IWL<9371> A_IWL<9370> A_IWL<9369> A_IWL<9368> A_IWL<9367> A_IWL<9366> A_IWL<9365> A_IWL<9364> A_IWL<9363> A_IWL<9362> A_IWL<9361> A_IWL<9360> A_IWL<9359> A_IWL<9358> A_IWL<9357> A_IWL<9356> A_IWL<9355> A_IWL<9354> A_IWL<9353> A_IWL<9352> A_IWL<9351> A_IWL<9350> A_IWL<9349> A_IWL<9348> A_IWL<9347> A_IWL<9346> A_IWL<9345> A_IWL<9344> A_IWL<9343> A_IWL<9342> A_IWL<9341> A_IWL<9340> A_IWL<9339> A_IWL<9338> A_IWL<9337> A_IWL<9336> A_IWL<9335> A_IWL<9334> A_IWL<9333> A_IWL<9332> A_IWL<9331> A_IWL<9330> A_IWL<9329> A_IWL<9328> A_IWL<9327> A_IWL<9326> A_IWL<9325> A_IWL<9324> A_IWL<9323> A_IWL<9322> A_IWL<9321> A_IWL<9320> A_IWL<9319> A_IWL<9318> A_IWL<9317> A_IWL<9316> A_IWL<9315> A_IWL<9314> A_IWL<9313> A_IWL<9312> A_IWL<9311> A_IWL<9310> A_IWL<9309> A_IWL<9308> A_IWL<9307> A_IWL<9306> A_IWL<9305> A_IWL<9304> A_IWL<9303> A_IWL<9302> A_IWL<9301> A_IWL<9300> A_IWL<9299> A_IWL<9298> A_IWL<9297> A_IWL<9296> A_IWL<9295> A_IWL<9294> A_IWL<9293> A_IWL<9292> A_IWL<9291> A_IWL<9290> A_IWL<9289> A_IWL<9288> A_IWL<9287> A_IWL<9286> A_IWL<9285> A_IWL<9284> A_IWL<9283> A_IWL<9282> A_IWL<9281> A_IWL<9280> A_IWL<9279> A_IWL<9278> A_IWL<9277> A_IWL<9276> A_IWL<9275> A_IWL<9274> A_IWL<9273> A_IWL<9272> A_IWL<9271> A_IWL<9270> A_IWL<9269> A_IWL<9268> A_IWL<9267> A_IWL<9266> A_IWL<9265> A_IWL<9264> A_IWL<9263> A_IWL<9262> A_IWL<9261> A_IWL<9260> A_IWL<9259> A_IWL<9258> A_IWL<9257> A_IWL<9256> A_IWL<9255> A_IWL<9254> A_IWL<9253> A_IWL<9252> A_IWL<9251> A_IWL<9250> A_IWL<9249> A_IWL<9248> A_IWL<9247> A_IWL<9246> A_IWL<9245> A_IWL<9244> A_IWL<9243> A_IWL<9242> A_IWL<9241> A_IWL<9240> A_IWL<9239> A_IWL<9238> A_IWL<9237> A_IWL<9236> A_IWL<9235> A_IWL<9234> A_IWL<9233> A_IWL<9232> A_IWL<9231> A_IWL<9230> A_IWL<9229> A_IWL<9228> A_IWL<9227> A_IWL<9226> A_IWL<9225> A_IWL<9224> A_IWL<9223> A_IWL<9222> A_IWL<9221> A_IWL<9220> A_IWL<9219> A_IWL<9218> A_IWL<9217> A_IWL<9216> A_IWL<10239> A_IWL<10238> A_IWL<10237> A_IWL<10236> A_IWL<10235> A_IWL<10234> A_IWL<10233> A_IWL<10232> A_IWL<10231> A_IWL<10230> A_IWL<10229> A_IWL<10228> A_IWL<10227> A_IWL<10226> A_IWL<10225> A_IWL<10224> A_IWL<10223> A_IWL<10222> A_IWL<10221> A_IWL<10220> A_IWL<10219> A_IWL<10218> A_IWL<10217> A_IWL<10216> A_IWL<10215> A_IWL<10214> A_IWL<10213> A_IWL<10212> A_IWL<10211> A_IWL<10210> A_IWL<10209> A_IWL<10208> A_IWL<10207> A_IWL<10206> A_IWL<10205> A_IWL<10204> A_IWL<10203> A_IWL<10202> A_IWL<10201> A_IWL<10200> A_IWL<10199> A_IWL<10198> A_IWL<10197> A_IWL<10196> A_IWL<10195> A_IWL<10194> A_IWL<10193> A_IWL<10192> A_IWL<10191> A_IWL<10190> A_IWL<10189> A_IWL<10188> A_IWL<10187> A_IWL<10186> A_IWL<10185> A_IWL<10184> A_IWL<10183> A_IWL<10182> A_IWL<10181> A_IWL<10180> A_IWL<10179> A_IWL<10178> A_IWL<10177> A_IWL<10176> A_IWL<10175> A_IWL<10174> A_IWL<10173> A_IWL<10172> A_IWL<10171> A_IWL<10170> A_IWL<10169> A_IWL<10168> A_IWL<10167> A_IWL<10166> A_IWL<10165> A_IWL<10164> A_IWL<10163> A_IWL<10162> A_IWL<10161> A_IWL<10160> A_IWL<10159> A_IWL<10158> A_IWL<10157> A_IWL<10156> A_IWL<10155> A_IWL<10154> A_IWL<10153> A_IWL<10152> A_IWL<10151> A_IWL<10150> A_IWL<10149> A_IWL<10148> A_IWL<10147> A_IWL<10146> A_IWL<10145> A_IWL<10144> A_IWL<10143> A_IWL<10142> A_IWL<10141> A_IWL<10140> A_IWL<10139> A_IWL<10138> A_IWL<10137> A_IWL<10136> A_IWL<10135> A_IWL<10134> A_IWL<10133> A_IWL<10132> A_IWL<10131> A_IWL<10130> A_IWL<10129> A_IWL<10128> A_IWL<10127> A_IWL<10126> A_IWL<10125> A_IWL<10124> A_IWL<10123> A_IWL<10122> A_IWL<10121> A_IWL<10120> A_IWL<10119> A_IWL<10118> A_IWL<10117> A_IWL<10116> A_IWL<10115> A_IWL<10114> A_IWL<10113> A_IWL<10112> A_IWL<10111> A_IWL<10110> A_IWL<10109> A_IWL<10108> A_IWL<10107> A_IWL<10106> A_IWL<10105> A_IWL<10104> A_IWL<10103> A_IWL<10102> A_IWL<10101> A_IWL<10100> A_IWL<10099> A_IWL<10098> A_IWL<10097> A_IWL<10096> A_IWL<10095> A_IWL<10094> A_IWL<10093> A_IWL<10092> A_IWL<10091> A_IWL<10090> A_IWL<10089> A_IWL<10088> A_IWL<10087> A_IWL<10086> A_IWL<10085> A_IWL<10084> A_IWL<10083> A_IWL<10082> A_IWL<10081> A_IWL<10080> A_IWL<10079> A_IWL<10078> A_IWL<10077> A_IWL<10076> A_IWL<10075> A_IWL<10074> A_IWL<10073> A_IWL<10072> A_IWL<10071> A_IWL<10070> A_IWL<10069> A_IWL<10068> A_IWL<10067> A_IWL<10066> A_IWL<10065> A_IWL<10064> A_IWL<10063> A_IWL<10062> A_IWL<10061> A_IWL<10060> A_IWL<10059> A_IWL<10058> A_IWL<10057> A_IWL<10056> A_IWL<10055> A_IWL<10054> A_IWL<10053> A_IWL<10052> A_IWL<10051> A_IWL<10050> A_IWL<10049> A_IWL<10048> A_IWL<10047> A_IWL<10046> A_IWL<10045> A_IWL<10044> A_IWL<10043> A_IWL<10042> A_IWL<10041> A_IWL<10040> A_IWL<10039> A_IWL<10038> A_IWL<10037> A_IWL<10036> A_IWL<10035> A_IWL<10034> A_IWL<10033> A_IWL<10032> A_IWL<10031> A_IWL<10030> A_IWL<10029> A_IWL<10028> A_IWL<10027> A_IWL<10026> A_IWL<10025> A_IWL<10024> A_IWL<10023> A_IWL<10022> A_IWL<10021> A_IWL<10020> A_IWL<10019> A_IWL<10018> A_IWL<10017> A_IWL<10016> A_IWL<10015> A_IWL<10014> A_IWL<10013> A_IWL<10012> A_IWL<10011> A_IWL<10010> A_IWL<10009> A_IWL<10008> A_IWL<10007> A_IWL<10006> A_IWL<10005> A_IWL<10004> A_IWL<10003> A_IWL<10002> A_IWL<10001> A_IWL<10000> A_IWL<9999> A_IWL<9998> A_IWL<9997> A_IWL<9996> A_IWL<9995> A_IWL<9994> A_IWL<9993> A_IWL<9992> A_IWL<9991> A_IWL<9990> A_IWL<9989> A_IWL<9988> A_IWL<9987> A_IWL<9986> A_IWL<9985> A_IWL<9984> A_IWL<9983> A_IWL<9982> A_IWL<9981> A_IWL<9980> A_IWL<9979> A_IWL<9978> A_IWL<9977> A_IWL<9976> A_IWL<9975> A_IWL<9974> A_IWL<9973> A_IWL<9972> A_IWL<9971> A_IWL<9970> A_IWL<9969> A_IWL<9968> A_IWL<9967> A_IWL<9966> A_IWL<9965> A_IWL<9964> A_IWL<9963> A_IWL<9962> A_IWL<9961> A_IWL<9960> A_IWL<9959> A_IWL<9958> A_IWL<9957> A_IWL<9956> A_IWL<9955> A_IWL<9954> A_IWL<9953> A_IWL<9952> A_IWL<9951> A_IWL<9950> A_IWL<9949> A_IWL<9948> A_IWL<9947> A_IWL<9946> A_IWL<9945> A_IWL<9944> A_IWL<9943> A_IWL<9942> A_IWL<9941> A_IWL<9940> A_IWL<9939> A_IWL<9938> A_IWL<9937> A_IWL<9936> A_IWL<9935> A_IWL<9934> A_IWL<9933> A_IWL<9932> A_IWL<9931> A_IWL<9930> A_IWL<9929> A_IWL<9928> A_IWL<9927> A_IWL<9926> A_IWL<9925> A_IWL<9924> A_IWL<9923> A_IWL<9922> A_IWL<9921> A_IWL<9920> A_IWL<9919> A_IWL<9918> A_IWL<9917> A_IWL<9916> A_IWL<9915> A_IWL<9914> A_IWL<9913> A_IWL<9912> A_IWL<9911> A_IWL<9910> A_IWL<9909> A_IWL<9908> A_IWL<9907> A_IWL<9906> A_IWL<9905> A_IWL<9904> A_IWL<9903> A_IWL<9902> A_IWL<9901> A_IWL<9900> A_IWL<9899> A_IWL<9898> A_IWL<9897> A_IWL<9896> A_IWL<9895> A_IWL<9894> A_IWL<9893> A_IWL<9892> A_IWL<9891> A_IWL<9890> A_IWL<9889> A_IWL<9888> A_IWL<9887> A_IWL<9886> A_IWL<9885> A_IWL<9884> A_IWL<9883> A_IWL<9882> A_IWL<9881> A_IWL<9880> A_IWL<9879> A_IWL<9878> A_IWL<9877> A_IWL<9876> A_IWL<9875> A_IWL<9874> A_IWL<9873> A_IWL<9872> A_IWL<9871> A_IWL<9870> A_IWL<9869> A_IWL<9868> A_IWL<9867> A_IWL<9866> A_IWL<9865> A_IWL<9864> A_IWL<9863> A_IWL<9862> A_IWL<9861> A_IWL<9860> A_IWL<9859> A_IWL<9858> A_IWL<9857> A_IWL<9856> A_IWL<9855> A_IWL<9854> A_IWL<9853> A_IWL<9852> A_IWL<9851> A_IWL<9850> A_IWL<9849> A_IWL<9848> A_IWL<9847> A_IWL<9846> A_IWL<9845> A_IWL<9844> A_IWL<9843> A_IWL<9842> A_IWL<9841> A_IWL<9840> A_IWL<9839> A_IWL<9838> A_IWL<9837> A_IWL<9836> A_IWL<9835> A_IWL<9834> A_IWL<9833> A_IWL<9832> A_IWL<9831> A_IWL<9830> A_IWL<9829> A_IWL<9828> A_IWL<9827> A_IWL<9826> A_IWL<9825> A_IWL<9824> A_IWL<9823> A_IWL<9822> A_IWL<9821> A_IWL<9820> A_IWL<9819> A_IWL<9818> A_IWL<9817> A_IWL<9816> A_IWL<9815> A_IWL<9814> A_IWL<9813> A_IWL<9812> A_IWL<9811> A_IWL<9810> A_IWL<9809> A_IWL<9808> A_IWL<9807> A_IWL<9806> A_IWL<9805> A_IWL<9804> A_IWL<9803> A_IWL<9802> A_IWL<9801> A_IWL<9800> A_IWL<9799> A_IWL<9798> A_IWL<9797> A_IWL<9796> A_IWL<9795> A_IWL<9794> A_IWL<9793> A_IWL<9792> A_IWL<9791> A_IWL<9790> A_IWL<9789> A_IWL<9788> A_IWL<9787> A_IWL<9786> A_IWL<9785> A_IWL<9784> A_IWL<9783> A_IWL<9782> A_IWL<9781> A_IWL<9780> A_IWL<9779> A_IWL<9778> A_IWL<9777> A_IWL<9776> A_IWL<9775> A_IWL<9774> A_IWL<9773> A_IWL<9772> A_IWL<9771> A_IWL<9770> A_IWL<9769> A_IWL<9768> A_IWL<9767> A_IWL<9766> A_IWL<9765> A_IWL<9764> A_IWL<9763> A_IWL<9762> A_IWL<9761> A_IWL<9760> A_IWL<9759> A_IWL<9758> A_IWL<9757> A_IWL<9756> A_IWL<9755> A_IWL<9754> A_IWL<9753> A_IWL<9752> A_IWL<9751> A_IWL<9750> A_IWL<9749> A_IWL<9748> A_IWL<9747> A_IWL<9746> A_IWL<9745> A_IWL<9744> A_IWL<9743> A_IWL<9742> A_IWL<9741> A_IWL<9740> A_IWL<9739> A_IWL<9738> A_IWL<9737> A_IWL<9736> A_IWL<9735> A_IWL<9734> A_IWL<9733> A_IWL<9732> A_IWL<9731> A_IWL<9730> A_IWL<9729> A_IWL<9728> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<18> A_BLC<37> A_BLC<36> A_BLC_TOP<37> A_BLC_TOP<36> A_BLT<37> A_BLT<36> A_BLT_TOP<37> A_BLT_TOP<36> A_IWL<9215> A_IWL<9214> A_IWL<9213> A_IWL<9212> A_IWL<9211> A_IWL<9210> A_IWL<9209> A_IWL<9208> A_IWL<9207> A_IWL<9206> A_IWL<9205> A_IWL<9204> A_IWL<9203> A_IWL<9202> A_IWL<9201> A_IWL<9200> A_IWL<9199> A_IWL<9198> A_IWL<9197> A_IWL<9196> A_IWL<9195> A_IWL<9194> A_IWL<9193> A_IWL<9192> A_IWL<9191> A_IWL<9190> A_IWL<9189> A_IWL<9188> A_IWL<9187> A_IWL<9186> A_IWL<9185> A_IWL<9184> A_IWL<9183> A_IWL<9182> A_IWL<9181> A_IWL<9180> A_IWL<9179> A_IWL<9178> A_IWL<9177> A_IWL<9176> A_IWL<9175> A_IWL<9174> A_IWL<9173> A_IWL<9172> A_IWL<9171> A_IWL<9170> A_IWL<9169> A_IWL<9168> A_IWL<9167> A_IWL<9166> A_IWL<9165> A_IWL<9164> A_IWL<9163> A_IWL<9162> A_IWL<9161> A_IWL<9160> A_IWL<9159> A_IWL<9158> A_IWL<9157> A_IWL<9156> A_IWL<9155> A_IWL<9154> A_IWL<9153> A_IWL<9152> A_IWL<9151> A_IWL<9150> A_IWL<9149> A_IWL<9148> A_IWL<9147> A_IWL<9146> A_IWL<9145> A_IWL<9144> A_IWL<9143> A_IWL<9142> A_IWL<9141> A_IWL<9140> A_IWL<9139> A_IWL<9138> A_IWL<9137> A_IWL<9136> A_IWL<9135> A_IWL<9134> A_IWL<9133> A_IWL<9132> A_IWL<9131> A_IWL<9130> A_IWL<9129> A_IWL<9128> A_IWL<9127> A_IWL<9126> A_IWL<9125> A_IWL<9124> A_IWL<9123> A_IWL<9122> A_IWL<9121> A_IWL<9120> A_IWL<9119> A_IWL<9118> A_IWL<9117> A_IWL<9116> A_IWL<9115> A_IWL<9114> A_IWL<9113> A_IWL<9112> A_IWL<9111> A_IWL<9110> A_IWL<9109> A_IWL<9108> A_IWL<9107> A_IWL<9106> A_IWL<9105> A_IWL<9104> A_IWL<9103> A_IWL<9102> A_IWL<9101> A_IWL<9100> A_IWL<9099> A_IWL<9098> A_IWL<9097> A_IWL<9096> A_IWL<9095> A_IWL<9094> A_IWL<9093> A_IWL<9092> A_IWL<9091> A_IWL<9090> A_IWL<9089> A_IWL<9088> A_IWL<9087> A_IWL<9086> A_IWL<9085> A_IWL<9084> A_IWL<9083> A_IWL<9082> A_IWL<9081> A_IWL<9080> A_IWL<9079> A_IWL<9078> A_IWL<9077> A_IWL<9076> A_IWL<9075> A_IWL<9074> A_IWL<9073> A_IWL<9072> A_IWL<9071> A_IWL<9070> A_IWL<9069> A_IWL<9068> A_IWL<9067> A_IWL<9066> A_IWL<9065> A_IWL<9064> A_IWL<9063> A_IWL<9062> A_IWL<9061> A_IWL<9060> A_IWL<9059> A_IWL<9058> A_IWL<9057> A_IWL<9056> A_IWL<9055> A_IWL<9054> A_IWL<9053> A_IWL<9052> A_IWL<9051> A_IWL<9050> A_IWL<9049> A_IWL<9048> A_IWL<9047> A_IWL<9046> A_IWL<9045> A_IWL<9044> A_IWL<9043> A_IWL<9042> A_IWL<9041> A_IWL<9040> A_IWL<9039> A_IWL<9038> A_IWL<9037> A_IWL<9036> A_IWL<9035> A_IWL<9034> A_IWL<9033> A_IWL<9032> A_IWL<9031> A_IWL<9030> A_IWL<9029> A_IWL<9028> A_IWL<9027> A_IWL<9026> A_IWL<9025> A_IWL<9024> A_IWL<9023> A_IWL<9022> A_IWL<9021> A_IWL<9020> A_IWL<9019> A_IWL<9018> A_IWL<9017> A_IWL<9016> A_IWL<9015> A_IWL<9014> A_IWL<9013> A_IWL<9012> A_IWL<9011> A_IWL<9010> A_IWL<9009> A_IWL<9008> A_IWL<9007> A_IWL<9006> A_IWL<9005> A_IWL<9004> A_IWL<9003> A_IWL<9002> A_IWL<9001> A_IWL<9000> A_IWL<8999> A_IWL<8998> A_IWL<8997> A_IWL<8996> A_IWL<8995> A_IWL<8994> A_IWL<8993> A_IWL<8992> A_IWL<8991> A_IWL<8990> A_IWL<8989> A_IWL<8988> A_IWL<8987> A_IWL<8986> A_IWL<8985> A_IWL<8984> A_IWL<8983> A_IWL<8982> A_IWL<8981> A_IWL<8980> A_IWL<8979> A_IWL<8978> A_IWL<8977> A_IWL<8976> A_IWL<8975> A_IWL<8974> A_IWL<8973> A_IWL<8972> A_IWL<8971> A_IWL<8970> A_IWL<8969> A_IWL<8968> A_IWL<8967> A_IWL<8966> A_IWL<8965> A_IWL<8964> A_IWL<8963> A_IWL<8962> A_IWL<8961> A_IWL<8960> A_IWL<8959> A_IWL<8958> A_IWL<8957> A_IWL<8956> A_IWL<8955> A_IWL<8954> A_IWL<8953> A_IWL<8952> A_IWL<8951> A_IWL<8950> A_IWL<8949> A_IWL<8948> A_IWL<8947> A_IWL<8946> A_IWL<8945> A_IWL<8944> A_IWL<8943> A_IWL<8942> A_IWL<8941> A_IWL<8940> A_IWL<8939> A_IWL<8938> A_IWL<8937> A_IWL<8936> A_IWL<8935> A_IWL<8934> A_IWL<8933> A_IWL<8932> A_IWL<8931> A_IWL<8930> A_IWL<8929> A_IWL<8928> A_IWL<8927> A_IWL<8926> A_IWL<8925> A_IWL<8924> A_IWL<8923> A_IWL<8922> A_IWL<8921> A_IWL<8920> A_IWL<8919> A_IWL<8918> A_IWL<8917> A_IWL<8916> A_IWL<8915> A_IWL<8914> A_IWL<8913> A_IWL<8912> A_IWL<8911> A_IWL<8910> A_IWL<8909> A_IWL<8908> A_IWL<8907> A_IWL<8906> A_IWL<8905> A_IWL<8904> A_IWL<8903> A_IWL<8902> A_IWL<8901> A_IWL<8900> A_IWL<8899> A_IWL<8898> A_IWL<8897> A_IWL<8896> A_IWL<8895> A_IWL<8894> A_IWL<8893> A_IWL<8892> A_IWL<8891> A_IWL<8890> A_IWL<8889> A_IWL<8888> A_IWL<8887> A_IWL<8886> A_IWL<8885> A_IWL<8884> A_IWL<8883> A_IWL<8882> A_IWL<8881> A_IWL<8880> A_IWL<8879> A_IWL<8878> A_IWL<8877> A_IWL<8876> A_IWL<8875> A_IWL<8874> A_IWL<8873> A_IWL<8872> A_IWL<8871> A_IWL<8870> A_IWL<8869> A_IWL<8868> A_IWL<8867> A_IWL<8866> A_IWL<8865> A_IWL<8864> A_IWL<8863> A_IWL<8862> A_IWL<8861> A_IWL<8860> A_IWL<8859> A_IWL<8858> A_IWL<8857> A_IWL<8856> A_IWL<8855> A_IWL<8854> A_IWL<8853> A_IWL<8852> A_IWL<8851> A_IWL<8850> A_IWL<8849> A_IWL<8848> A_IWL<8847> A_IWL<8846> A_IWL<8845> A_IWL<8844> A_IWL<8843> A_IWL<8842> A_IWL<8841> A_IWL<8840> A_IWL<8839> A_IWL<8838> A_IWL<8837> A_IWL<8836> A_IWL<8835> A_IWL<8834> A_IWL<8833> A_IWL<8832> A_IWL<8831> A_IWL<8830> A_IWL<8829> A_IWL<8828> A_IWL<8827> A_IWL<8826> A_IWL<8825> A_IWL<8824> A_IWL<8823> A_IWL<8822> A_IWL<8821> A_IWL<8820> A_IWL<8819> A_IWL<8818> A_IWL<8817> A_IWL<8816> A_IWL<8815> A_IWL<8814> A_IWL<8813> A_IWL<8812> A_IWL<8811> A_IWL<8810> A_IWL<8809> A_IWL<8808> A_IWL<8807> A_IWL<8806> A_IWL<8805> A_IWL<8804> A_IWL<8803> A_IWL<8802> A_IWL<8801> A_IWL<8800> A_IWL<8799> A_IWL<8798> A_IWL<8797> A_IWL<8796> A_IWL<8795> A_IWL<8794> A_IWL<8793> A_IWL<8792> A_IWL<8791> A_IWL<8790> A_IWL<8789> A_IWL<8788> A_IWL<8787> A_IWL<8786> A_IWL<8785> A_IWL<8784> A_IWL<8783> A_IWL<8782> A_IWL<8781> A_IWL<8780> A_IWL<8779> A_IWL<8778> A_IWL<8777> A_IWL<8776> A_IWL<8775> A_IWL<8774> A_IWL<8773> A_IWL<8772> A_IWL<8771> A_IWL<8770> A_IWL<8769> A_IWL<8768> A_IWL<8767> A_IWL<8766> A_IWL<8765> A_IWL<8764> A_IWL<8763> A_IWL<8762> A_IWL<8761> A_IWL<8760> A_IWL<8759> A_IWL<8758> A_IWL<8757> A_IWL<8756> A_IWL<8755> A_IWL<8754> A_IWL<8753> A_IWL<8752> A_IWL<8751> A_IWL<8750> A_IWL<8749> A_IWL<8748> A_IWL<8747> A_IWL<8746> A_IWL<8745> A_IWL<8744> A_IWL<8743> A_IWL<8742> A_IWL<8741> A_IWL<8740> A_IWL<8739> A_IWL<8738> A_IWL<8737> A_IWL<8736> A_IWL<8735> A_IWL<8734> A_IWL<8733> A_IWL<8732> A_IWL<8731> A_IWL<8730> A_IWL<8729> A_IWL<8728> A_IWL<8727> A_IWL<8726> A_IWL<8725> A_IWL<8724> A_IWL<8723> A_IWL<8722> A_IWL<8721> A_IWL<8720> A_IWL<8719> A_IWL<8718> A_IWL<8717> A_IWL<8716> A_IWL<8715> A_IWL<8714> A_IWL<8713> A_IWL<8712> A_IWL<8711> A_IWL<8710> A_IWL<8709> A_IWL<8708> A_IWL<8707> A_IWL<8706> A_IWL<8705> A_IWL<8704> A_IWL<9727> A_IWL<9726> A_IWL<9725> A_IWL<9724> A_IWL<9723> A_IWL<9722> A_IWL<9721> A_IWL<9720> A_IWL<9719> A_IWL<9718> A_IWL<9717> A_IWL<9716> A_IWL<9715> A_IWL<9714> A_IWL<9713> A_IWL<9712> A_IWL<9711> A_IWL<9710> A_IWL<9709> A_IWL<9708> A_IWL<9707> A_IWL<9706> A_IWL<9705> A_IWL<9704> A_IWL<9703> A_IWL<9702> A_IWL<9701> A_IWL<9700> A_IWL<9699> A_IWL<9698> A_IWL<9697> A_IWL<9696> A_IWL<9695> A_IWL<9694> A_IWL<9693> A_IWL<9692> A_IWL<9691> A_IWL<9690> A_IWL<9689> A_IWL<9688> A_IWL<9687> A_IWL<9686> A_IWL<9685> A_IWL<9684> A_IWL<9683> A_IWL<9682> A_IWL<9681> A_IWL<9680> A_IWL<9679> A_IWL<9678> A_IWL<9677> A_IWL<9676> A_IWL<9675> A_IWL<9674> A_IWL<9673> A_IWL<9672> A_IWL<9671> A_IWL<9670> A_IWL<9669> A_IWL<9668> A_IWL<9667> A_IWL<9666> A_IWL<9665> A_IWL<9664> A_IWL<9663> A_IWL<9662> A_IWL<9661> A_IWL<9660> A_IWL<9659> A_IWL<9658> A_IWL<9657> A_IWL<9656> A_IWL<9655> A_IWL<9654> A_IWL<9653> A_IWL<9652> A_IWL<9651> A_IWL<9650> A_IWL<9649> A_IWL<9648> A_IWL<9647> A_IWL<9646> A_IWL<9645> A_IWL<9644> A_IWL<9643> A_IWL<9642> A_IWL<9641> A_IWL<9640> A_IWL<9639> A_IWL<9638> A_IWL<9637> A_IWL<9636> A_IWL<9635> A_IWL<9634> A_IWL<9633> A_IWL<9632> A_IWL<9631> A_IWL<9630> A_IWL<9629> A_IWL<9628> A_IWL<9627> A_IWL<9626> A_IWL<9625> A_IWL<9624> A_IWL<9623> A_IWL<9622> A_IWL<9621> A_IWL<9620> A_IWL<9619> A_IWL<9618> A_IWL<9617> A_IWL<9616> A_IWL<9615> A_IWL<9614> A_IWL<9613> A_IWL<9612> A_IWL<9611> A_IWL<9610> A_IWL<9609> A_IWL<9608> A_IWL<9607> A_IWL<9606> A_IWL<9605> A_IWL<9604> A_IWL<9603> A_IWL<9602> A_IWL<9601> A_IWL<9600> A_IWL<9599> A_IWL<9598> A_IWL<9597> A_IWL<9596> A_IWL<9595> A_IWL<9594> A_IWL<9593> A_IWL<9592> A_IWL<9591> A_IWL<9590> A_IWL<9589> A_IWL<9588> A_IWL<9587> A_IWL<9586> A_IWL<9585> A_IWL<9584> A_IWL<9583> A_IWL<9582> A_IWL<9581> A_IWL<9580> A_IWL<9579> A_IWL<9578> A_IWL<9577> A_IWL<9576> A_IWL<9575> A_IWL<9574> A_IWL<9573> A_IWL<9572> A_IWL<9571> A_IWL<9570> A_IWL<9569> A_IWL<9568> A_IWL<9567> A_IWL<9566> A_IWL<9565> A_IWL<9564> A_IWL<9563> A_IWL<9562> A_IWL<9561> A_IWL<9560> A_IWL<9559> A_IWL<9558> A_IWL<9557> A_IWL<9556> A_IWL<9555> A_IWL<9554> A_IWL<9553> A_IWL<9552> A_IWL<9551> A_IWL<9550> A_IWL<9549> A_IWL<9548> A_IWL<9547> A_IWL<9546> A_IWL<9545> A_IWL<9544> A_IWL<9543> A_IWL<9542> A_IWL<9541> A_IWL<9540> A_IWL<9539> A_IWL<9538> A_IWL<9537> A_IWL<9536> A_IWL<9535> A_IWL<9534> A_IWL<9533> A_IWL<9532> A_IWL<9531> A_IWL<9530> A_IWL<9529> A_IWL<9528> A_IWL<9527> A_IWL<9526> A_IWL<9525> A_IWL<9524> A_IWL<9523> A_IWL<9522> A_IWL<9521> A_IWL<9520> A_IWL<9519> A_IWL<9518> A_IWL<9517> A_IWL<9516> A_IWL<9515> A_IWL<9514> A_IWL<9513> A_IWL<9512> A_IWL<9511> A_IWL<9510> A_IWL<9509> A_IWL<9508> A_IWL<9507> A_IWL<9506> A_IWL<9505> A_IWL<9504> A_IWL<9503> A_IWL<9502> A_IWL<9501> A_IWL<9500> A_IWL<9499> A_IWL<9498> A_IWL<9497> A_IWL<9496> A_IWL<9495> A_IWL<9494> A_IWL<9493> A_IWL<9492> A_IWL<9491> A_IWL<9490> A_IWL<9489> A_IWL<9488> A_IWL<9487> A_IWL<9486> A_IWL<9485> A_IWL<9484> A_IWL<9483> A_IWL<9482> A_IWL<9481> A_IWL<9480> A_IWL<9479> A_IWL<9478> A_IWL<9477> A_IWL<9476> A_IWL<9475> A_IWL<9474> A_IWL<9473> A_IWL<9472> A_IWL<9471> A_IWL<9470> A_IWL<9469> A_IWL<9468> A_IWL<9467> A_IWL<9466> A_IWL<9465> A_IWL<9464> A_IWL<9463> A_IWL<9462> A_IWL<9461> A_IWL<9460> A_IWL<9459> A_IWL<9458> A_IWL<9457> A_IWL<9456> A_IWL<9455> A_IWL<9454> A_IWL<9453> A_IWL<9452> A_IWL<9451> A_IWL<9450> A_IWL<9449> A_IWL<9448> A_IWL<9447> A_IWL<9446> A_IWL<9445> A_IWL<9444> A_IWL<9443> A_IWL<9442> A_IWL<9441> A_IWL<9440> A_IWL<9439> A_IWL<9438> A_IWL<9437> A_IWL<9436> A_IWL<9435> A_IWL<9434> A_IWL<9433> A_IWL<9432> A_IWL<9431> A_IWL<9430> A_IWL<9429> A_IWL<9428> A_IWL<9427> A_IWL<9426> A_IWL<9425> A_IWL<9424> A_IWL<9423> A_IWL<9422> A_IWL<9421> A_IWL<9420> A_IWL<9419> A_IWL<9418> A_IWL<9417> A_IWL<9416> A_IWL<9415> A_IWL<9414> A_IWL<9413> A_IWL<9412> A_IWL<9411> A_IWL<9410> A_IWL<9409> A_IWL<9408> A_IWL<9407> A_IWL<9406> A_IWL<9405> A_IWL<9404> A_IWL<9403> A_IWL<9402> A_IWL<9401> A_IWL<9400> A_IWL<9399> A_IWL<9398> A_IWL<9397> A_IWL<9396> A_IWL<9395> A_IWL<9394> A_IWL<9393> A_IWL<9392> A_IWL<9391> A_IWL<9390> A_IWL<9389> A_IWL<9388> A_IWL<9387> A_IWL<9386> A_IWL<9385> A_IWL<9384> A_IWL<9383> A_IWL<9382> A_IWL<9381> A_IWL<9380> A_IWL<9379> A_IWL<9378> A_IWL<9377> A_IWL<9376> A_IWL<9375> A_IWL<9374> A_IWL<9373> A_IWL<9372> A_IWL<9371> A_IWL<9370> A_IWL<9369> A_IWL<9368> A_IWL<9367> A_IWL<9366> A_IWL<9365> A_IWL<9364> A_IWL<9363> A_IWL<9362> A_IWL<9361> A_IWL<9360> A_IWL<9359> A_IWL<9358> A_IWL<9357> A_IWL<9356> A_IWL<9355> A_IWL<9354> A_IWL<9353> A_IWL<9352> A_IWL<9351> A_IWL<9350> A_IWL<9349> A_IWL<9348> A_IWL<9347> A_IWL<9346> A_IWL<9345> A_IWL<9344> A_IWL<9343> A_IWL<9342> A_IWL<9341> A_IWL<9340> A_IWL<9339> A_IWL<9338> A_IWL<9337> A_IWL<9336> A_IWL<9335> A_IWL<9334> A_IWL<9333> A_IWL<9332> A_IWL<9331> A_IWL<9330> A_IWL<9329> A_IWL<9328> A_IWL<9327> A_IWL<9326> A_IWL<9325> A_IWL<9324> A_IWL<9323> A_IWL<9322> A_IWL<9321> A_IWL<9320> A_IWL<9319> A_IWL<9318> A_IWL<9317> A_IWL<9316> A_IWL<9315> A_IWL<9314> A_IWL<9313> A_IWL<9312> A_IWL<9311> A_IWL<9310> A_IWL<9309> A_IWL<9308> A_IWL<9307> A_IWL<9306> A_IWL<9305> A_IWL<9304> A_IWL<9303> A_IWL<9302> A_IWL<9301> A_IWL<9300> A_IWL<9299> A_IWL<9298> A_IWL<9297> A_IWL<9296> A_IWL<9295> A_IWL<9294> A_IWL<9293> A_IWL<9292> A_IWL<9291> A_IWL<9290> A_IWL<9289> A_IWL<9288> A_IWL<9287> A_IWL<9286> A_IWL<9285> A_IWL<9284> A_IWL<9283> A_IWL<9282> A_IWL<9281> A_IWL<9280> A_IWL<9279> A_IWL<9278> A_IWL<9277> A_IWL<9276> A_IWL<9275> A_IWL<9274> A_IWL<9273> A_IWL<9272> A_IWL<9271> A_IWL<9270> A_IWL<9269> A_IWL<9268> A_IWL<9267> A_IWL<9266> A_IWL<9265> A_IWL<9264> A_IWL<9263> A_IWL<9262> A_IWL<9261> A_IWL<9260> A_IWL<9259> A_IWL<9258> A_IWL<9257> A_IWL<9256> A_IWL<9255> A_IWL<9254> A_IWL<9253> A_IWL<9252> A_IWL<9251> A_IWL<9250> A_IWL<9249> A_IWL<9248> A_IWL<9247> A_IWL<9246> A_IWL<9245> A_IWL<9244> A_IWL<9243> A_IWL<9242> A_IWL<9241> A_IWL<9240> A_IWL<9239> A_IWL<9238> A_IWL<9237> A_IWL<9236> A_IWL<9235> A_IWL<9234> A_IWL<9233> A_IWL<9232> A_IWL<9231> A_IWL<9230> A_IWL<9229> A_IWL<9228> A_IWL<9227> A_IWL<9226> A_IWL<9225> A_IWL<9224> A_IWL<9223> A_IWL<9222> A_IWL<9221> A_IWL<9220> A_IWL<9219> A_IWL<9218> A_IWL<9217> A_IWL<9216> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<17> A_BLC<35> A_BLC<34> A_BLC_TOP<35> A_BLC_TOP<34> A_BLT<35> A_BLT<34> A_BLT_TOP<35> A_BLT_TOP<34> A_IWL<8703> A_IWL<8702> A_IWL<8701> A_IWL<8700> A_IWL<8699> A_IWL<8698> A_IWL<8697> A_IWL<8696> A_IWL<8695> A_IWL<8694> A_IWL<8693> A_IWL<8692> A_IWL<8691> A_IWL<8690> A_IWL<8689> A_IWL<8688> A_IWL<8687> A_IWL<8686> A_IWL<8685> A_IWL<8684> A_IWL<8683> A_IWL<8682> A_IWL<8681> A_IWL<8680> A_IWL<8679> A_IWL<8678> A_IWL<8677> A_IWL<8676> A_IWL<8675> A_IWL<8674> A_IWL<8673> A_IWL<8672> A_IWL<8671> A_IWL<8670> A_IWL<8669> A_IWL<8668> A_IWL<8667> A_IWL<8666> A_IWL<8665> A_IWL<8664> A_IWL<8663> A_IWL<8662> A_IWL<8661> A_IWL<8660> A_IWL<8659> A_IWL<8658> A_IWL<8657> A_IWL<8656> A_IWL<8655> A_IWL<8654> A_IWL<8653> A_IWL<8652> A_IWL<8651> A_IWL<8650> A_IWL<8649> A_IWL<8648> A_IWL<8647> A_IWL<8646> A_IWL<8645> A_IWL<8644> A_IWL<8643> A_IWL<8642> A_IWL<8641> A_IWL<8640> A_IWL<8639> A_IWL<8638> A_IWL<8637> A_IWL<8636> A_IWL<8635> A_IWL<8634> A_IWL<8633> A_IWL<8632> A_IWL<8631> A_IWL<8630> A_IWL<8629> A_IWL<8628> A_IWL<8627> A_IWL<8626> A_IWL<8625> A_IWL<8624> A_IWL<8623> A_IWL<8622> A_IWL<8621> A_IWL<8620> A_IWL<8619> A_IWL<8618> A_IWL<8617> A_IWL<8616> A_IWL<8615> A_IWL<8614> A_IWL<8613> A_IWL<8612> A_IWL<8611> A_IWL<8610> A_IWL<8609> A_IWL<8608> A_IWL<8607> A_IWL<8606> A_IWL<8605> A_IWL<8604> A_IWL<8603> A_IWL<8602> A_IWL<8601> A_IWL<8600> A_IWL<8599> A_IWL<8598> A_IWL<8597> A_IWL<8596> A_IWL<8595> A_IWL<8594> A_IWL<8593> A_IWL<8592> A_IWL<8591> A_IWL<8590> A_IWL<8589> A_IWL<8588> A_IWL<8587> A_IWL<8586> A_IWL<8585> A_IWL<8584> A_IWL<8583> A_IWL<8582> A_IWL<8581> A_IWL<8580> A_IWL<8579> A_IWL<8578> A_IWL<8577> A_IWL<8576> A_IWL<8575> A_IWL<8574> A_IWL<8573> A_IWL<8572> A_IWL<8571> A_IWL<8570> A_IWL<8569> A_IWL<8568> A_IWL<8567> A_IWL<8566> A_IWL<8565> A_IWL<8564> A_IWL<8563> A_IWL<8562> A_IWL<8561> A_IWL<8560> A_IWL<8559> A_IWL<8558> A_IWL<8557> A_IWL<8556> A_IWL<8555> A_IWL<8554> A_IWL<8553> A_IWL<8552> A_IWL<8551> A_IWL<8550> A_IWL<8549> A_IWL<8548> A_IWL<8547> A_IWL<8546> A_IWL<8545> A_IWL<8544> A_IWL<8543> A_IWL<8542> A_IWL<8541> A_IWL<8540> A_IWL<8539> A_IWL<8538> A_IWL<8537> A_IWL<8536> A_IWL<8535> A_IWL<8534> A_IWL<8533> A_IWL<8532> A_IWL<8531> A_IWL<8530> A_IWL<8529> A_IWL<8528> A_IWL<8527> A_IWL<8526> A_IWL<8525> A_IWL<8524> A_IWL<8523> A_IWL<8522> A_IWL<8521> A_IWL<8520> A_IWL<8519> A_IWL<8518> A_IWL<8517> A_IWL<8516> A_IWL<8515> A_IWL<8514> A_IWL<8513> A_IWL<8512> A_IWL<8511> A_IWL<8510> A_IWL<8509> A_IWL<8508> A_IWL<8507> A_IWL<8506> A_IWL<8505> A_IWL<8504> A_IWL<8503> A_IWL<8502> A_IWL<8501> A_IWL<8500> A_IWL<8499> A_IWL<8498> A_IWL<8497> A_IWL<8496> A_IWL<8495> A_IWL<8494> A_IWL<8493> A_IWL<8492> A_IWL<8491> A_IWL<8490> A_IWL<8489> A_IWL<8488> A_IWL<8487> A_IWL<8486> A_IWL<8485> A_IWL<8484> A_IWL<8483> A_IWL<8482> A_IWL<8481> A_IWL<8480> A_IWL<8479> A_IWL<8478> A_IWL<8477> A_IWL<8476> A_IWL<8475> A_IWL<8474> A_IWL<8473> A_IWL<8472> A_IWL<8471> A_IWL<8470> A_IWL<8469> A_IWL<8468> A_IWL<8467> A_IWL<8466> A_IWL<8465> A_IWL<8464> A_IWL<8463> A_IWL<8462> A_IWL<8461> A_IWL<8460> A_IWL<8459> A_IWL<8458> A_IWL<8457> A_IWL<8456> A_IWL<8455> A_IWL<8454> A_IWL<8453> A_IWL<8452> A_IWL<8451> A_IWL<8450> A_IWL<8449> A_IWL<8448> A_IWL<8447> A_IWL<8446> A_IWL<8445> A_IWL<8444> A_IWL<8443> A_IWL<8442> A_IWL<8441> A_IWL<8440> A_IWL<8439> A_IWL<8438> A_IWL<8437> A_IWL<8436> A_IWL<8435> A_IWL<8434> A_IWL<8433> A_IWL<8432> A_IWL<8431> A_IWL<8430> A_IWL<8429> A_IWL<8428> A_IWL<8427> A_IWL<8426> A_IWL<8425> A_IWL<8424> A_IWL<8423> A_IWL<8422> A_IWL<8421> A_IWL<8420> A_IWL<8419> A_IWL<8418> A_IWL<8417> A_IWL<8416> A_IWL<8415> A_IWL<8414> A_IWL<8413> A_IWL<8412> A_IWL<8411> A_IWL<8410> A_IWL<8409> A_IWL<8408> A_IWL<8407> A_IWL<8406> A_IWL<8405> A_IWL<8404> A_IWL<8403> A_IWL<8402> A_IWL<8401> A_IWL<8400> A_IWL<8399> A_IWL<8398> A_IWL<8397> A_IWL<8396> A_IWL<8395> A_IWL<8394> A_IWL<8393> A_IWL<8392> A_IWL<8391> A_IWL<8390> A_IWL<8389> A_IWL<8388> A_IWL<8387> A_IWL<8386> A_IWL<8385> A_IWL<8384> A_IWL<8383> A_IWL<8382> A_IWL<8381> A_IWL<8380> A_IWL<8379> A_IWL<8378> A_IWL<8377> A_IWL<8376> A_IWL<8375> A_IWL<8374> A_IWL<8373> A_IWL<8372> A_IWL<8371> A_IWL<8370> A_IWL<8369> A_IWL<8368> A_IWL<8367> A_IWL<8366> A_IWL<8365> A_IWL<8364> A_IWL<8363> A_IWL<8362> A_IWL<8361> A_IWL<8360> A_IWL<8359> A_IWL<8358> A_IWL<8357> A_IWL<8356> A_IWL<8355> A_IWL<8354> A_IWL<8353> A_IWL<8352> A_IWL<8351> A_IWL<8350> A_IWL<8349> A_IWL<8348> A_IWL<8347> A_IWL<8346> A_IWL<8345> A_IWL<8344> A_IWL<8343> A_IWL<8342> A_IWL<8341> A_IWL<8340> A_IWL<8339> A_IWL<8338> A_IWL<8337> A_IWL<8336> A_IWL<8335> A_IWL<8334> A_IWL<8333> A_IWL<8332> A_IWL<8331> A_IWL<8330> A_IWL<8329> A_IWL<8328> A_IWL<8327> A_IWL<8326> A_IWL<8325> A_IWL<8324> A_IWL<8323> A_IWL<8322> A_IWL<8321> A_IWL<8320> A_IWL<8319> A_IWL<8318> A_IWL<8317> A_IWL<8316> A_IWL<8315> A_IWL<8314> A_IWL<8313> A_IWL<8312> A_IWL<8311> A_IWL<8310> A_IWL<8309> A_IWL<8308> A_IWL<8307> A_IWL<8306> A_IWL<8305> A_IWL<8304> A_IWL<8303> A_IWL<8302> A_IWL<8301> A_IWL<8300> A_IWL<8299> A_IWL<8298> A_IWL<8297> A_IWL<8296> A_IWL<8295> A_IWL<8294> A_IWL<8293> A_IWL<8292> A_IWL<8291> A_IWL<8290> A_IWL<8289> A_IWL<8288> A_IWL<8287> A_IWL<8286> A_IWL<8285> A_IWL<8284> A_IWL<8283> A_IWL<8282> A_IWL<8281> A_IWL<8280> A_IWL<8279> A_IWL<8278> A_IWL<8277> A_IWL<8276> A_IWL<8275> A_IWL<8274> A_IWL<8273> A_IWL<8272> A_IWL<8271> A_IWL<8270> A_IWL<8269> A_IWL<8268> A_IWL<8267> A_IWL<8266> A_IWL<8265> A_IWL<8264> A_IWL<8263> A_IWL<8262> A_IWL<8261> A_IWL<8260> A_IWL<8259> A_IWL<8258> A_IWL<8257> A_IWL<8256> A_IWL<8255> A_IWL<8254> A_IWL<8253> A_IWL<8252> A_IWL<8251> A_IWL<8250> A_IWL<8249> A_IWL<8248> A_IWL<8247> A_IWL<8246> A_IWL<8245> A_IWL<8244> A_IWL<8243> A_IWL<8242> A_IWL<8241> A_IWL<8240> A_IWL<8239> A_IWL<8238> A_IWL<8237> A_IWL<8236> A_IWL<8235> A_IWL<8234> A_IWL<8233> A_IWL<8232> A_IWL<8231> A_IWL<8230> A_IWL<8229> A_IWL<8228> A_IWL<8227> A_IWL<8226> A_IWL<8225> A_IWL<8224> A_IWL<8223> A_IWL<8222> A_IWL<8221> A_IWL<8220> A_IWL<8219> A_IWL<8218> A_IWL<8217> A_IWL<8216> A_IWL<8215> A_IWL<8214> A_IWL<8213> A_IWL<8212> A_IWL<8211> A_IWL<8210> A_IWL<8209> A_IWL<8208> A_IWL<8207> A_IWL<8206> A_IWL<8205> A_IWL<8204> A_IWL<8203> A_IWL<8202> A_IWL<8201> A_IWL<8200> A_IWL<8199> A_IWL<8198> A_IWL<8197> A_IWL<8196> A_IWL<8195> A_IWL<8194> A_IWL<8193> A_IWL<8192> A_IWL<9215> A_IWL<9214> A_IWL<9213> A_IWL<9212> A_IWL<9211> A_IWL<9210> A_IWL<9209> A_IWL<9208> A_IWL<9207> A_IWL<9206> A_IWL<9205> A_IWL<9204> A_IWL<9203> A_IWL<9202> A_IWL<9201> A_IWL<9200> A_IWL<9199> A_IWL<9198> A_IWL<9197> A_IWL<9196> A_IWL<9195> A_IWL<9194> A_IWL<9193> A_IWL<9192> A_IWL<9191> A_IWL<9190> A_IWL<9189> A_IWL<9188> A_IWL<9187> A_IWL<9186> A_IWL<9185> A_IWL<9184> A_IWL<9183> A_IWL<9182> A_IWL<9181> A_IWL<9180> A_IWL<9179> A_IWL<9178> A_IWL<9177> A_IWL<9176> A_IWL<9175> A_IWL<9174> A_IWL<9173> A_IWL<9172> A_IWL<9171> A_IWL<9170> A_IWL<9169> A_IWL<9168> A_IWL<9167> A_IWL<9166> A_IWL<9165> A_IWL<9164> A_IWL<9163> A_IWL<9162> A_IWL<9161> A_IWL<9160> A_IWL<9159> A_IWL<9158> A_IWL<9157> A_IWL<9156> A_IWL<9155> A_IWL<9154> A_IWL<9153> A_IWL<9152> A_IWL<9151> A_IWL<9150> A_IWL<9149> A_IWL<9148> A_IWL<9147> A_IWL<9146> A_IWL<9145> A_IWL<9144> A_IWL<9143> A_IWL<9142> A_IWL<9141> A_IWL<9140> A_IWL<9139> A_IWL<9138> A_IWL<9137> A_IWL<9136> A_IWL<9135> A_IWL<9134> A_IWL<9133> A_IWL<9132> A_IWL<9131> A_IWL<9130> A_IWL<9129> A_IWL<9128> A_IWL<9127> A_IWL<9126> A_IWL<9125> A_IWL<9124> A_IWL<9123> A_IWL<9122> A_IWL<9121> A_IWL<9120> A_IWL<9119> A_IWL<9118> A_IWL<9117> A_IWL<9116> A_IWL<9115> A_IWL<9114> A_IWL<9113> A_IWL<9112> A_IWL<9111> A_IWL<9110> A_IWL<9109> A_IWL<9108> A_IWL<9107> A_IWL<9106> A_IWL<9105> A_IWL<9104> A_IWL<9103> A_IWL<9102> A_IWL<9101> A_IWL<9100> A_IWL<9099> A_IWL<9098> A_IWL<9097> A_IWL<9096> A_IWL<9095> A_IWL<9094> A_IWL<9093> A_IWL<9092> A_IWL<9091> A_IWL<9090> A_IWL<9089> A_IWL<9088> A_IWL<9087> A_IWL<9086> A_IWL<9085> A_IWL<9084> A_IWL<9083> A_IWL<9082> A_IWL<9081> A_IWL<9080> A_IWL<9079> A_IWL<9078> A_IWL<9077> A_IWL<9076> A_IWL<9075> A_IWL<9074> A_IWL<9073> A_IWL<9072> A_IWL<9071> A_IWL<9070> A_IWL<9069> A_IWL<9068> A_IWL<9067> A_IWL<9066> A_IWL<9065> A_IWL<9064> A_IWL<9063> A_IWL<9062> A_IWL<9061> A_IWL<9060> A_IWL<9059> A_IWL<9058> A_IWL<9057> A_IWL<9056> A_IWL<9055> A_IWL<9054> A_IWL<9053> A_IWL<9052> A_IWL<9051> A_IWL<9050> A_IWL<9049> A_IWL<9048> A_IWL<9047> A_IWL<9046> A_IWL<9045> A_IWL<9044> A_IWL<9043> A_IWL<9042> A_IWL<9041> A_IWL<9040> A_IWL<9039> A_IWL<9038> A_IWL<9037> A_IWL<9036> A_IWL<9035> A_IWL<9034> A_IWL<9033> A_IWL<9032> A_IWL<9031> A_IWL<9030> A_IWL<9029> A_IWL<9028> A_IWL<9027> A_IWL<9026> A_IWL<9025> A_IWL<9024> A_IWL<9023> A_IWL<9022> A_IWL<9021> A_IWL<9020> A_IWL<9019> A_IWL<9018> A_IWL<9017> A_IWL<9016> A_IWL<9015> A_IWL<9014> A_IWL<9013> A_IWL<9012> A_IWL<9011> A_IWL<9010> A_IWL<9009> A_IWL<9008> A_IWL<9007> A_IWL<9006> A_IWL<9005> A_IWL<9004> A_IWL<9003> A_IWL<9002> A_IWL<9001> A_IWL<9000> A_IWL<8999> A_IWL<8998> A_IWL<8997> A_IWL<8996> A_IWL<8995> A_IWL<8994> A_IWL<8993> A_IWL<8992> A_IWL<8991> A_IWL<8990> A_IWL<8989> A_IWL<8988> A_IWL<8987> A_IWL<8986> A_IWL<8985> A_IWL<8984> A_IWL<8983> A_IWL<8982> A_IWL<8981> A_IWL<8980> A_IWL<8979> A_IWL<8978> A_IWL<8977> A_IWL<8976> A_IWL<8975> A_IWL<8974> A_IWL<8973> A_IWL<8972> A_IWL<8971> A_IWL<8970> A_IWL<8969> A_IWL<8968> A_IWL<8967> A_IWL<8966> A_IWL<8965> A_IWL<8964> A_IWL<8963> A_IWL<8962> A_IWL<8961> A_IWL<8960> A_IWL<8959> A_IWL<8958> A_IWL<8957> A_IWL<8956> A_IWL<8955> A_IWL<8954> A_IWL<8953> A_IWL<8952> A_IWL<8951> A_IWL<8950> A_IWL<8949> A_IWL<8948> A_IWL<8947> A_IWL<8946> A_IWL<8945> A_IWL<8944> A_IWL<8943> A_IWL<8942> A_IWL<8941> A_IWL<8940> A_IWL<8939> A_IWL<8938> A_IWL<8937> A_IWL<8936> A_IWL<8935> A_IWL<8934> A_IWL<8933> A_IWL<8932> A_IWL<8931> A_IWL<8930> A_IWL<8929> A_IWL<8928> A_IWL<8927> A_IWL<8926> A_IWL<8925> A_IWL<8924> A_IWL<8923> A_IWL<8922> A_IWL<8921> A_IWL<8920> A_IWL<8919> A_IWL<8918> A_IWL<8917> A_IWL<8916> A_IWL<8915> A_IWL<8914> A_IWL<8913> A_IWL<8912> A_IWL<8911> A_IWL<8910> A_IWL<8909> A_IWL<8908> A_IWL<8907> A_IWL<8906> A_IWL<8905> A_IWL<8904> A_IWL<8903> A_IWL<8902> A_IWL<8901> A_IWL<8900> A_IWL<8899> A_IWL<8898> A_IWL<8897> A_IWL<8896> A_IWL<8895> A_IWL<8894> A_IWL<8893> A_IWL<8892> A_IWL<8891> A_IWL<8890> A_IWL<8889> A_IWL<8888> A_IWL<8887> A_IWL<8886> A_IWL<8885> A_IWL<8884> A_IWL<8883> A_IWL<8882> A_IWL<8881> A_IWL<8880> A_IWL<8879> A_IWL<8878> A_IWL<8877> A_IWL<8876> A_IWL<8875> A_IWL<8874> A_IWL<8873> A_IWL<8872> A_IWL<8871> A_IWL<8870> A_IWL<8869> A_IWL<8868> A_IWL<8867> A_IWL<8866> A_IWL<8865> A_IWL<8864> A_IWL<8863> A_IWL<8862> A_IWL<8861> A_IWL<8860> A_IWL<8859> A_IWL<8858> A_IWL<8857> A_IWL<8856> A_IWL<8855> A_IWL<8854> A_IWL<8853> A_IWL<8852> A_IWL<8851> A_IWL<8850> A_IWL<8849> A_IWL<8848> A_IWL<8847> A_IWL<8846> A_IWL<8845> A_IWL<8844> A_IWL<8843> A_IWL<8842> A_IWL<8841> A_IWL<8840> A_IWL<8839> A_IWL<8838> A_IWL<8837> A_IWL<8836> A_IWL<8835> A_IWL<8834> A_IWL<8833> A_IWL<8832> A_IWL<8831> A_IWL<8830> A_IWL<8829> A_IWL<8828> A_IWL<8827> A_IWL<8826> A_IWL<8825> A_IWL<8824> A_IWL<8823> A_IWL<8822> A_IWL<8821> A_IWL<8820> A_IWL<8819> A_IWL<8818> A_IWL<8817> A_IWL<8816> A_IWL<8815> A_IWL<8814> A_IWL<8813> A_IWL<8812> A_IWL<8811> A_IWL<8810> A_IWL<8809> A_IWL<8808> A_IWL<8807> A_IWL<8806> A_IWL<8805> A_IWL<8804> A_IWL<8803> A_IWL<8802> A_IWL<8801> A_IWL<8800> A_IWL<8799> A_IWL<8798> A_IWL<8797> A_IWL<8796> A_IWL<8795> A_IWL<8794> A_IWL<8793> A_IWL<8792> A_IWL<8791> A_IWL<8790> A_IWL<8789> A_IWL<8788> A_IWL<8787> A_IWL<8786> A_IWL<8785> A_IWL<8784> A_IWL<8783> A_IWL<8782> A_IWL<8781> A_IWL<8780> A_IWL<8779> A_IWL<8778> A_IWL<8777> A_IWL<8776> A_IWL<8775> A_IWL<8774> A_IWL<8773> A_IWL<8772> A_IWL<8771> A_IWL<8770> A_IWL<8769> A_IWL<8768> A_IWL<8767> A_IWL<8766> A_IWL<8765> A_IWL<8764> A_IWL<8763> A_IWL<8762> A_IWL<8761> A_IWL<8760> A_IWL<8759> A_IWL<8758> A_IWL<8757> A_IWL<8756> A_IWL<8755> A_IWL<8754> A_IWL<8753> A_IWL<8752> A_IWL<8751> A_IWL<8750> A_IWL<8749> A_IWL<8748> A_IWL<8747> A_IWL<8746> A_IWL<8745> A_IWL<8744> A_IWL<8743> A_IWL<8742> A_IWL<8741> A_IWL<8740> A_IWL<8739> A_IWL<8738> A_IWL<8737> A_IWL<8736> A_IWL<8735> A_IWL<8734> A_IWL<8733> A_IWL<8732> A_IWL<8731> A_IWL<8730> A_IWL<8729> A_IWL<8728> A_IWL<8727> A_IWL<8726> A_IWL<8725> A_IWL<8724> A_IWL<8723> A_IWL<8722> A_IWL<8721> A_IWL<8720> A_IWL<8719> A_IWL<8718> A_IWL<8717> A_IWL<8716> A_IWL<8715> A_IWL<8714> A_IWL<8713> A_IWL<8712> A_IWL<8711> A_IWL<8710> A_IWL<8709> A_IWL<8708> A_IWL<8707> A_IWL<8706> A_IWL<8705> A_IWL<8704> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<16> A_BLC<33> A_BLC<32> A_BLC_TOP<33> A_BLC_TOP<32> A_BLT<33> A_BLT<32> A_BLT_TOP<33> A_BLT_TOP<32> A_IWL<8191> A_IWL<8190> A_IWL<8189> A_IWL<8188> A_IWL<8187> A_IWL<8186> A_IWL<8185> A_IWL<8184> A_IWL<8183> A_IWL<8182> A_IWL<8181> A_IWL<8180> A_IWL<8179> A_IWL<8178> A_IWL<8177> A_IWL<8176> A_IWL<8175> A_IWL<8174> A_IWL<8173> A_IWL<8172> A_IWL<8171> A_IWL<8170> A_IWL<8169> A_IWL<8168> A_IWL<8167> A_IWL<8166> A_IWL<8165> A_IWL<8164> A_IWL<8163> A_IWL<8162> A_IWL<8161> A_IWL<8160> A_IWL<8159> A_IWL<8158> A_IWL<8157> A_IWL<8156> A_IWL<8155> A_IWL<8154> A_IWL<8153> A_IWL<8152> A_IWL<8151> A_IWL<8150> A_IWL<8149> A_IWL<8148> A_IWL<8147> A_IWL<8146> A_IWL<8145> A_IWL<8144> A_IWL<8143> A_IWL<8142> A_IWL<8141> A_IWL<8140> A_IWL<8139> A_IWL<8138> A_IWL<8137> A_IWL<8136> A_IWL<8135> A_IWL<8134> A_IWL<8133> A_IWL<8132> A_IWL<8131> A_IWL<8130> A_IWL<8129> A_IWL<8128> A_IWL<8127> A_IWL<8126> A_IWL<8125> A_IWL<8124> A_IWL<8123> A_IWL<8122> A_IWL<8121> A_IWL<8120> A_IWL<8119> A_IWL<8118> A_IWL<8117> A_IWL<8116> A_IWL<8115> A_IWL<8114> A_IWL<8113> A_IWL<8112> A_IWL<8111> A_IWL<8110> A_IWL<8109> A_IWL<8108> A_IWL<8107> A_IWL<8106> A_IWL<8105> A_IWL<8104> A_IWL<8103> A_IWL<8102> A_IWL<8101> A_IWL<8100> A_IWL<8099> A_IWL<8098> A_IWL<8097> A_IWL<8096> A_IWL<8095> A_IWL<8094> A_IWL<8093> A_IWL<8092> A_IWL<8091> A_IWL<8090> A_IWL<8089> A_IWL<8088> A_IWL<8087> A_IWL<8086> A_IWL<8085> A_IWL<8084> A_IWL<8083> A_IWL<8082> A_IWL<8081> A_IWL<8080> A_IWL<8079> A_IWL<8078> A_IWL<8077> A_IWL<8076> A_IWL<8075> A_IWL<8074> A_IWL<8073> A_IWL<8072> A_IWL<8071> A_IWL<8070> A_IWL<8069> A_IWL<8068> A_IWL<8067> A_IWL<8066> A_IWL<8065> A_IWL<8064> A_IWL<8063> A_IWL<8062> A_IWL<8061> A_IWL<8060> A_IWL<8059> A_IWL<8058> A_IWL<8057> A_IWL<8056> A_IWL<8055> A_IWL<8054> A_IWL<8053> A_IWL<8052> A_IWL<8051> A_IWL<8050> A_IWL<8049> A_IWL<8048> A_IWL<8047> A_IWL<8046> A_IWL<8045> A_IWL<8044> A_IWL<8043> A_IWL<8042> A_IWL<8041> A_IWL<8040> A_IWL<8039> A_IWL<8038> A_IWL<8037> A_IWL<8036> A_IWL<8035> A_IWL<8034> A_IWL<8033> A_IWL<8032> A_IWL<8031> A_IWL<8030> A_IWL<8029> A_IWL<8028> A_IWL<8027> A_IWL<8026> A_IWL<8025> A_IWL<8024> A_IWL<8023> A_IWL<8022> A_IWL<8021> A_IWL<8020> A_IWL<8019> A_IWL<8018> A_IWL<8017> A_IWL<8016> A_IWL<8015> A_IWL<8014> A_IWL<8013> A_IWL<8012> A_IWL<8011> A_IWL<8010> A_IWL<8009> A_IWL<8008> A_IWL<8007> A_IWL<8006> A_IWL<8005> A_IWL<8004> A_IWL<8003> A_IWL<8002> A_IWL<8001> A_IWL<8000> A_IWL<7999> A_IWL<7998> A_IWL<7997> A_IWL<7996> A_IWL<7995> A_IWL<7994> A_IWL<7993> A_IWL<7992> A_IWL<7991> A_IWL<7990> A_IWL<7989> A_IWL<7988> A_IWL<7987> A_IWL<7986> A_IWL<7985> A_IWL<7984> A_IWL<7983> A_IWL<7982> A_IWL<7981> A_IWL<7980> A_IWL<7979> A_IWL<7978> A_IWL<7977> A_IWL<7976> A_IWL<7975> A_IWL<7974> A_IWL<7973> A_IWL<7972> A_IWL<7971> A_IWL<7970> A_IWL<7969> A_IWL<7968> A_IWL<7967> A_IWL<7966> A_IWL<7965> A_IWL<7964> A_IWL<7963> A_IWL<7962> A_IWL<7961> A_IWL<7960> A_IWL<7959> A_IWL<7958> A_IWL<7957> A_IWL<7956> A_IWL<7955> A_IWL<7954> A_IWL<7953> A_IWL<7952> A_IWL<7951> A_IWL<7950> A_IWL<7949> A_IWL<7948> A_IWL<7947> A_IWL<7946> A_IWL<7945> A_IWL<7944> A_IWL<7943> A_IWL<7942> A_IWL<7941> A_IWL<7940> A_IWL<7939> A_IWL<7938> A_IWL<7937> A_IWL<7936> A_IWL<7935> A_IWL<7934> A_IWL<7933> A_IWL<7932> A_IWL<7931> A_IWL<7930> A_IWL<7929> A_IWL<7928> A_IWL<7927> A_IWL<7926> A_IWL<7925> A_IWL<7924> A_IWL<7923> A_IWL<7922> A_IWL<7921> A_IWL<7920> A_IWL<7919> A_IWL<7918> A_IWL<7917> A_IWL<7916> A_IWL<7915> A_IWL<7914> A_IWL<7913> A_IWL<7912> A_IWL<7911> A_IWL<7910> A_IWL<7909> A_IWL<7908> A_IWL<7907> A_IWL<7906> A_IWL<7905> A_IWL<7904> A_IWL<7903> A_IWL<7902> A_IWL<7901> A_IWL<7900> A_IWL<7899> A_IWL<7898> A_IWL<7897> A_IWL<7896> A_IWL<7895> A_IWL<7894> A_IWL<7893> A_IWL<7892> A_IWL<7891> A_IWL<7890> A_IWL<7889> A_IWL<7888> A_IWL<7887> A_IWL<7886> A_IWL<7885> A_IWL<7884> A_IWL<7883> A_IWL<7882> A_IWL<7881> A_IWL<7880> A_IWL<7879> A_IWL<7878> A_IWL<7877> A_IWL<7876> A_IWL<7875> A_IWL<7874> A_IWL<7873> A_IWL<7872> A_IWL<7871> A_IWL<7870> A_IWL<7869> A_IWL<7868> A_IWL<7867> A_IWL<7866> A_IWL<7865> A_IWL<7864> A_IWL<7863> A_IWL<7862> A_IWL<7861> A_IWL<7860> A_IWL<7859> A_IWL<7858> A_IWL<7857> A_IWL<7856> A_IWL<7855> A_IWL<7854> A_IWL<7853> A_IWL<7852> A_IWL<7851> A_IWL<7850> A_IWL<7849> A_IWL<7848> A_IWL<7847> A_IWL<7846> A_IWL<7845> A_IWL<7844> A_IWL<7843> A_IWL<7842> A_IWL<7841> A_IWL<7840> A_IWL<7839> A_IWL<7838> A_IWL<7837> A_IWL<7836> A_IWL<7835> A_IWL<7834> A_IWL<7833> A_IWL<7832> A_IWL<7831> A_IWL<7830> A_IWL<7829> A_IWL<7828> A_IWL<7827> A_IWL<7826> A_IWL<7825> A_IWL<7824> A_IWL<7823> A_IWL<7822> A_IWL<7821> A_IWL<7820> A_IWL<7819> A_IWL<7818> A_IWL<7817> A_IWL<7816> A_IWL<7815> A_IWL<7814> A_IWL<7813> A_IWL<7812> A_IWL<7811> A_IWL<7810> A_IWL<7809> A_IWL<7808> A_IWL<7807> A_IWL<7806> A_IWL<7805> A_IWL<7804> A_IWL<7803> A_IWL<7802> A_IWL<7801> A_IWL<7800> A_IWL<7799> A_IWL<7798> A_IWL<7797> A_IWL<7796> A_IWL<7795> A_IWL<7794> A_IWL<7793> A_IWL<7792> A_IWL<7791> A_IWL<7790> A_IWL<7789> A_IWL<7788> A_IWL<7787> A_IWL<7786> A_IWL<7785> A_IWL<7784> A_IWL<7783> A_IWL<7782> A_IWL<7781> A_IWL<7780> A_IWL<7779> A_IWL<7778> A_IWL<7777> A_IWL<7776> A_IWL<7775> A_IWL<7774> A_IWL<7773> A_IWL<7772> A_IWL<7771> A_IWL<7770> A_IWL<7769> A_IWL<7768> A_IWL<7767> A_IWL<7766> A_IWL<7765> A_IWL<7764> A_IWL<7763> A_IWL<7762> A_IWL<7761> A_IWL<7760> A_IWL<7759> A_IWL<7758> A_IWL<7757> A_IWL<7756> A_IWL<7755> A_IWL<7754> A_IWL<7753> A_IWL<7752> A_IWL<7751> A_IWL<7750> A_IWL<7749> A_IWL<7748> A_IWL<7747> A_IWL<7746> A_IWL<7745> A_IWL<7744> A_IWL<7743> A_IWL<7742> A_IWL<7741> A_IWL<7740> A_IWL<7739> A_IWL<7738> A_IWL<7737> A_IWL<7736> A_IWL<7735> A_IWL<7734> A_IWL<7733> A_IWL<7732> A_IWL<7731> A_IWL<7730> A_IWL<7729> A_IWL<7728> A_IWL<7727> A_IWL<7726> A_IWL<7725> A_IWL<7724> A_IWL<7723> A_IWL<7722> A_IWL<7721> A_IWL<7720> A_IWL<7719> A_IWL<7718> A_IWL<7717> A_IWL<7716> A_IWL<7715> A_IWL<7714> A_IWL<7713> A_IWL<7712> A_IWL<7711> A_IWL<7710> A_IWL<7709> A_IWL<7708> A_IWL<7707> A_IWL<7706> A_IWL<7705> A_IWL<7704> A_IWL<7703> A_IWL<7702> A_IWL<7701> A_IWL<7700> A_IWL<7699> A_IWL<7698> A_IWL<7697> A_IWL<7696> A_IWL<7695> A_IWL<7694> A_IWL<7693> A_IWL<7692> A_IWL<7691> A_IWL<7690> A_IWL<7689> A_IWL<7688> A_IWL<7687> A_IWL<7686> A_IWL<7685> A_IWL<7684> A_IWL<7683> A_IWL<7682> A_IWL<7681> A_IWL<7680> A_IWL<8703> A_IWL<8702> A_IWL<8701> A_IWL<8700> A_IWL<8699> A_IWL<8698> A_IWL<8697> A_IWL<8696> A_IWL<8695> A_IWL<8694> A_IWL<8693> A_IWL<8692> A_IWL<8691> A_IWL<8690> A_IWL<8689> A_IWL<8688> A_IWL<8687> A_IWL<8686> A_IWL<8685> A_IWL<8684> A_IWL<8683> A_IWL<8682> A_IWL<8681> A_IWL<8680> A_IWL<8679> A_IWL<8678> A_IWL<8677> A_IWL<8676> A_IWL<8675> A_IWL<8674> A_IWL<8673> A_IWL<8672> A_IWL<8671> A_IWL<8670> A_IWL<8669> A_IWL<8668> A_IWL<8667> A_IWL<8666> A_IWL<8665> A_IWL<8664> A_IWL<8663> A_IWL<8662> A_IWL<8661> A_IWL<8660> A_IWL<8659> A_IWL<8658> A_IWL<8657> A_IWL<8656> A_IWL<8655> A_IWL<8654> A_IWL<8653> A_IWL<8652> A_IWL<8651> A_IWL<8650> A_IWL<8649> A_IWL<8648> A_IWL<8647> A_IWL<8646> A_IWL<8645> A_IWL<8644> A_IWL<8643> A_IWL<8642> A_IWL<8641> A_IWL<8640> A_IWL<8639> A_IWL<8638> A_IWL<8637> A_IWL<8636> A_IWL<8635> A_IWL<8634> A_IWL<8633> A_IWL<8632> A_IWL<8631> A_IWL<8630> A_IWL<8629> A_IWL<8628> A_IWL<8627> A_IWL<8626> A_IWL<8625> A_IWL<8624> A_IWL<8623> A_IWL<8622> A_IWL<8621> A_IWL<8620> A_IWL<8619> A_IWL<8618> A_IWL<8617> A_IWL<8616> A_IWL<8615> A_IWL<8614> A_IWL<8613> A_IWL<8612> A_IWL<8611> A_IWL<8610> A_IWL<8609> A_IWL<8608> A_IWL<8607> A_IWL<8606> A_IWL<8605> A_IWL<8604> A_IWL<8603> A_IWL<8602> A_IWL<8601> A_IWL<8600> A_IWL<8599> A_IWL<8598> A_IWL<8597> A_IWL<8596> A_IWL<8595> A_IWL<8594> A_IWL<8593> A_IWL<8592> A_IWL<8591> A_IWL<8590> A_IWL<8589> A_IWL<8588> A_IWL<8587> A_IWL<8586> A_IWL<8585> A_IWL<8584> A_IWL<8583> A_IWL<8582> A_IWL<8581> A_IWL<8580> A_IWL<8579> A_IWL<8578> A_IWL<8577> A_IWL<8576> A_IWL<8575> A_IWL<8574> A_IWL<8573> A_IWL<8572> A_IWL<8571> A_IWL<8570> A_IWL<8569> A_IWL<8568> A_IWL<8567> A_IWL<8566> A_IWL<8565> A_IWL<8564> A_IWL<8563> A_IWL<8562> A_IWL<8561> A_IWL<8560> A_IWL<8559> A_IWL<8558> A_IWL<8557> A_IWL<8556> A_IWL<8555> A_IWL<8554> A_IWL<8553> A_IWL<8552> A_IWL<8551> A_IWL<8550> A_IWL<8549> A_IWL<8548> A_IWL<8547> A_IWL<8546> A_IWL<8545> A_IWL<8544> A_IWL<8543> A_IWL<8542> A_IWL<8541> A_IWL<8540> A_IWL<8539> A_IWL<8538> A_IWL<8537> A_IWL<8536> A_IWL<8535> A_IWL<8534> A_IWL<8533> A_IWL<8532> A_IWL<8531> A_IWL<8530> A_IWL<8529> A_IWL<8528> A_IWL<8527> A_IWL<8526> A_IWL<8525> A_IWL<8524> A_IWL<8523> A_IWL<8522> A_IWL<8521> A_IWL<8520> A_IWL<8519> A_IWL<8518> A_IWL<8517> A_IWL<8516> A_IWL<8515> A_IWL<8514> A_IWL<8513> A_IWL<8512> A_IWL<8511> A_IWL<8510> A_IWL<8509> A_IWL<8508> A_IWL<8507> A_IWL<8506> A_IWL<8505> A_IWL<8504> A_IWL<8503> A_IWL<8502> A_IWL<8501> A_IWL<8500> A_IWL<8499> A_IWL<8498> A_IWL<8497> A_IWL<8496> A_IWL<8495> A_IWL<8494> A_IWL<8493> A_IWL<8492> A_IWL<8491> A_IWL<8490> A_IWL<8489> A_IWL<8488> A_IWL<8487> A_IWL<8486> A_IWL<8485> A_IWL<8484> A_IWL<8483> A_IWL<8482> A_IWL<8481> A_IWL<8480> A_IWL<8479> A_IWL<8478> A_IWL<8477> A_IWL<8476> A_IWL<8475> A_IWL<8474> A_IWL<8473> A_IWL<8472> A_IWL<8471> A_IWL<8470> A_IWL<8469> A_IWL<8468> A_IWL<8467> A_IWL<8466> A_IWL<8465> A_IWL<8464> A_IWL<8463> A_IWL<8462> A_IWL<8461> A_IWL<8460> A_IWL<8459> A_IWL<8458> A_IWL<8457> A_IWL<8456> A_IWL<8455> A_IWL<8454> A_IWL<8453> A_IWL<8452> A_IWL<8451> A_IWL<8450> A_IWL<8449> A_IWL<8448> A_IWL<8447> A_IWL<8446> A_IWL<8445> A_IWL<8444> A_IWL<8443> A_IWL<8442> A_IWL<8441> A_IWL<8440> A_IWL<8439> A_IWL<8438> A_IWL<8437> A_IWL<8436> A_IWL<8435> A_IWL<8434> A_IWL<8433> A_IWL<8432> A_IWL<8431> A_IWL<8430> A_IWL<8429> A_IWL<8428> A_IWL<8427> A_IWL<8426> A_IWL<8425> A_IWL<8424> A_IWL<8423> A_IWL<8422> A_IWL<8421> A_IWL<8420> A_IWL<8419> A_IWL<8418> A_IWL<8417> A_IWL<8416> A_IWL<8415> A_IWL<8414> A_IWL<8413> A_IWL<8412> A_IWL<8411> A_IWL<8410> A_IWL<8409> A_IWL<8408> A_IWL<8407> A_IWL<8406> A_IWL<8405> A_IWL<8404> A_IWL<8403> A_IWL<8402> A_IWL<8401> A_IWL<8400> A_IWL<8399> A_IWL<8398> A_IWL<8397> A_IWL<8396> A_IWL<8395> A_IWL<8394> A_IWL<8393> A_IWL<8392> A_IWL<8391> A_IWL<8390> A_IWL<8389> A_IWL<8388> A_IWL<8387> A_IWL<8386> A_IWL<8385> A_IWL<8384> A_IWL<8383> A_IWL<8382> A_IWL<8381> A_IWL<8380> A_IWL<8379> A_IWL<8378> A_IWL<8377> A_IWL<8376> A_IWL<8375> A_IWL<8374> A_IWL<8373> A_IWL<8372> A_IWL<8371> A_IWL<8370> A_IWL<8369> A_IWL<8368> A_IWL<8367> A_IWL<8366> A_IWL<8365> A_IWL<8364> A_IWL<8363> A_IWL<8362> A_IWL<8361> A_IWL<8360> A_IWL<8359> A_IWL<8358> A_IWL<8357> A_IWL<8356> A_IWL<8355> A_IWL<8354> A_IWL<8353> A_IWL<8352> A_IWL<8351> A_IWL<8350> A_IWL<8349> A_IWL<8348> A_IWL<8347> A_IWL<8346> A_IWL<8345> A_IWL<8344> A_IWL<8343> A_IWL<8342> A_IWL<8341> A_IWL<8340> A_IWL<8339> A_IWL<8338> A_IWL<8337> A_IWL<8336> A_IWL<8335> A_IWL<8334> A_IWL<8333> A_IWL<8332> A_IWL<8331> A_IWL<8330> A_IWL<8329> A_IWL<8328> A_IWL<8327> A_IWL<8326> A_IWL<8325> A_IWL<8324> A_IWL<8323> A_IWL<8322> A_IWL<8321> A_IWL<8320> A_IWL<8319> A_IWL<8318> A_IWL<8317> A_IWL<8316> A_IWL<8315> A_IWL<8314> A_IWL<8313> A_IWL<8312> A_IWL<8311> A_IWL<8310> A_IWL<8309> A_IWL<8308> A_IWL<8307> A_IWL<8306> A_IWL<8305> A_IWL<8304> A_IWL<8303> A_IWL<8302> A_IWL<8301> A_IWL<8300> A_IWL<8299> A_IWL<8298> A_IWL<8297> A_IWL<8296> A_IWL<8295> A_IWL<8294> A_IWL<8293> A_IWL<8292> A_IWL<8291> A_IWL<8290> A_IWL<8289> A_IWL<8288> A_IWL<8287> A_IWL<8286> A_IWL<8285> A_IWL<8284> A_IWL<8283> A_IWL<8282> A_IWL<8281> A_IWL<8280> A_IWL<8279> A_IWL<8278> A_IWL<8277> A_IWL<8276> A_IWL<8275> A_IWL<8274> A_IWL<8273> A_IWL<8272> A_IWL<8271> A_IWL<8270> A_IWL<8269> A_IWL<8268> A_IWL<8267> A_IWL<8266> A_IWL<8265> A_IWL<8264> A_IWL<8263> A_IWL<8262> A_IWL<8261> A_IWL<8260> A_IWL<8259> A_IWL<8258> A_IWL<8257> A_IWL<8256> A_IWL<8255> A_IWL<8254> A_IWL<8253> A_IWL<8252> A_IWL<8251> A_IWL<8250> A_IWL<8249> A_IWL<8248> A_IWL<8247> A_IWL<8246> A_IWL<8245> A_IWL<8244> A_IWL<8243> A_IWL<8242> A_IWL<8241> A_IWL<8240> A_IWL<8239> A_IWL<8238> A_IWL<8237> A_IWL<8236> A_IWL<8235> A_IWL<8234> A_IWL<8233> A_IWL<8232> A_IWL<8231> A_IWL<8230> A_IWL<8229> A_IWL<8228> A_IWL<8227> A_IWL<8226> A_IWL<8225> A_IWL<8224> A_IWL<8223> A_IWL<8222> A_IWL<8221> A_IWL<8220> A_IWL<8219> A_IWL<8218> A_IWL<8217> A_IWL<8216> A_IWL<8215> A_IWL<8214> A_IWL<8213> A_IWL<8212> A_IWL<8211> A_IWL<8210> A_IWL<8209> A_IWL<8208> A_IWL<8207> A_IWL<8206> A_IWL<8205> A_IWL<8204> A_IWL<8203> A_IWL<8202> A_IWL<8201> A_IWL<8200> A_IWL<8199> A_IWL<8198> A_IWL<8197> A_IWL<8196> A_IWL<8195> A_IWL<8194> A_IWL<8193> A_IWL<8192> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<15> A_BLC<31> A_BLC<30> A_BLC_TOP<31> A_BLC_TOP<30> A_BLT<31> A_BLT<30> A_BLT_TOP<31> A_BLT_TOP<30> A_IWL<7679> A_IWL<7678> A_IWL<7677> A_IWL<7676> A_IWL<7675> A_IWL<7674> A_IWL<7673> A_IWL<7672> A_IWL<7671> A_IWL<7670> A_IWL<7669> A_IWL<7668> A_IWL<7667> A_IWL<7666> A_IWL<7665> A_IWL<7664> A_IWL<7663> A_IWL<7662> A_IWL<7661> A_IWL<7660> A_IWL<7659> A_IWL<7658> A_IWL<7657> A_IWL<7656> A_IWL<7655> A_IWL<7654> A_IWL<7653> A_IWL<7652> A_IWL<7651> A_IWL<7650> A_IWL<7649> A_IWL<7648> A_IWL<7647> A_IWL<7646> A_IWL<7645> A_IWL<7644> A_IWL<7643> A_IWL<7642> A_IWL<7641> A_IWL<7640> A_IWL<7639> A_IWL<7638> A_IWL<7637> A_IWL<7636> A_IWL<7635> A_IWL<7634> A_IWL<7633> A_IWL<7632> A_IWL<7631> A_IWL<7630> A_IWL<7629> A_IWL<7628> A_IWL<7627> A_IWL<7626> A_IWL<7625> A_IWL<7624> A_IWL<7623> A_IWL<7622> A_IWL<7621> A_IWL<7620> A_IWL<7619> A_IWL<7618> A_IWL<7617> A_IWL<7616> A_IWL<7615> A_IWL<7614> A_IWL<7613> A_IWL<7612> A_IWL<7611> A_IWL<7610> A_IWL<7609> A_IWL<7608> A_IWL<7607> A_IWL<7606> A_IWL<7605> A_IWL<7604> A_IWL<7603> A_IWL<7602> A_IWL<7601> A_IWL<7600> A_IWL<7599> A_IWL<7598> A_IWL<7597> A_IWL<7596> A_IWL<7595> A_IWL<7594> A_IWL<7593> A_IWL<7592> A_IWL<7591> A_IWL<7590> A_IWL<7589> A_IWL<7588> A_IWL<7587> A_IWL<7586> A_IWL<7585> A_IWL<7584> A_IWL<7583> A_IWL<7582> A_IWL<7581> A_IWL<7580> A_IWL<7579> A_IWL<7578> A_IWL<7577> A_IWL<7576> A_IWL<7575> A_IWL<7574> A_IWL<7573> A_IWL<7572> A_IWL<7571> A_IWL<7570> A_IWL<7569> A_IWL<7568> A_IWL<7567> A_IWL<7566> A_IWL<7565> A_IWL<7564> A_IWL<7563> A_IWL<7562> A_IWL<7561> A_IWL<7560> A_IWL<7559> A_IWL<7558> A_IWL<7557> A_IWL<7556> A_IWL<7555> A_IWL<7554> A_IWL<7553> A_IWL<7552> A_IWL<7551> A_IWL<7550> A_IWL<7549> A_IWL<7548> A_IWL<7547> A_IWL<7546> A_IWL<7545> A_IWL<7544> A_IWL<7543> A_IWL<7542> A_IWL<7541> A_IWL<7540> A_IWL<7539> A_IWL<7538> A_IWL<7537> A_IWL<7536> A_IWL<7535> A_IWL<7534> A_IWL<7533> A_IWL<7532> A_IWL<7531> A_IWL<7530> A_IWL<7529> A_IWL<7528> A_IWL<7527> A_IWL<7526> A_IWL<7525> A_IWL<7524> A_IWL<7523> A_IWL<7522> A_IWL<7521> A_IWL<7520> A_IWL<7519> A_IWL<7518> A_IWL<7517> A_IWL<7516> A_IWL<7515> A_IWL<7514> A_IWL<7513> A_IWL<7512> A_IWL<7511> A_IWL<7510> A_IWL<7509> A_IWL<7508> A_IWL<7507> A_IWL<7506> A_IWL<7505> A_IWL<7504> A_IWL<7503> A_IWL<7502> A_IWL<7501> A_IWL<7500> A_IWL<7499> A_IWL<7498> A_IWL<7497> A_IWL<7496> A_IWL<7495> A_IWL<7494> A_IWL<7493> A_IWL<7492> A_IWL<7491> A_IWL<7490> A_IWL<7489> A_IWL<7488> A_IWL<7487> A_IWL<7486> A_IWL<7485> A_IWL<7484> A_IWL<7483> A_IWL<7482> A_IWL<7481> A_IWL<7480> A_IWL<7479> A_IWL<7478> A_IWL<7477> A_IWL<7476> A_IWL<7475> A_IWL<7474> A_IWL<7473> A_IWL<7472> A_IWL<7471> A_IWL<7470> A_IWL<7469> A_IWL<7468> A_IWL<7467> A_IWL<7466> A_IWL<7465> A_IWL<7464> A_IWL<7463> A_IWL<7462> A_IWL<7461> A_IWL<7460> A_IWL<7459> A_IWL<7458> A_IWL<7457> A_IWL<7456> A_IWL<7455> A_IWL<7454> A_IWL<7453> A_IWL<7452> A_IWL<7451> A_IWL<7450> A_IWL<7449> A_IWL<7448> A_IWL<7447> A_IWL<7446> A_IWL<7445> A_IWL<7444> A_IWL<7443> A_IWL<7442> A_IWL<7441> A_IWL<7440> A_IWL<7439> A_IWL<7438> A_IWL<7437> A_IWL<7436> A_IWL<7435> A_IWL<7434> A_IWL<7433> A_IWL<7432> A_IWL<7431> A_IWL<7430> A_IWL<7429> A_IWL<7428> A_IWL<7427> A_IWL<7426> A_IWL<7425> A_IWL<7424> A_IWL<7423> A_IWL<7422> A_IWL<7421> A_IWL<7420> A_IWL<7419> A_IWL<7418> A_IWL<7417> A_IWL<7416> A_IWL<7415> A_IWL<7414> A_IWL<7413> A_IWL<7412> A_IWL<7411> A_IWL<7410> A_IWL<7409> A_IWL<7408> A_IWL<7407> A_IWL<7406> A_IWL<7405> A_IWL<7404> A_IWL<7403> A_IWL<7402> A_IWL<7401> A_IWL<7400> A_IWL<7399> A_IWL<7398> A_IWL<7397> A_IWL<7396> A_IWL<7395> A_IWL<7394> A_IWL<7393> A_IWL<7392> A_IWL<7391> A_IWL<7390> A_IWL<7389> A_IWL<7388> A_IWL<7387> A_IWL<7386> A_IWL<7385> A_IWL<7384> A_IWL<7383> A_IWL<7382> A_IWL<7381> A_IWL<7380> A_IWL<7379> A_IWL<7378> A_IWL<7377> A_IWL<7376> A_IWL<7375> A_IWL<7374> A_IWL<7373> A_IWL<7372> A_IWL<7371> A_IWL<7370> A_IWL<7369> A_IWL<7368> A_IWL<7367> A_IWL<7366> A_IWL<7365> A_IWL<7364> A_IWL<7363> A_IWL<7362> A_IWL<7361> A_IWL<7360> A_IWL<7359> A_IWL<7358> A_IWL<7357> A_IWL<7356> A_IWL<7355> A_IWL<7354> A_IWL<7353> A_IWL<7352> A_IWL<7351> A_IWL<7350> A_IWL<7349> A_IWL<7348> A_IWL<7347> A_IWL<7346> A_IWL<7345> A_IWL<7344> A_IWL<7343> A_IWL<7342> A_IWL<7341> A_IWL<7340> A_IWL<7339> A_IWL<7338> A_IWL<7337> A_IWL<7336> A_IWL<7335> A_IWL<7334> A_IWL<7333> A_IWL<7332> A_IWL<7331> A_IWL<7330> A_IWL<7329> A_IWL<7328> A_IWL<7327> A_IWL<7326> A_IWL<7325> A_IWL<7324> A_IWL<7323> A_IWL<7322> A_IWL<7321> A_IWL<7320> A_IWL<7319> A_IWL<7318> A_IWL<7317> A_IWL<7316> A_IWL<7315> A_IWL<7314> A_IWL<7313> A_IWL<7312> A_IWL<7311> A_IWL<7310> A_IWL<7309> A_IWL<7308> A_IWL<7307> A_IWL<7306> A_IWL<7305> A_IWL<7304> A_IWL<7303> A_IWL<7302> A_IWL<7301> A_IWL<7300> A_IWL<7299> A_IWL<7298> A_IWL<7297> A_IWL<7296> A_IWL<7295> A_IWL<7294> A_IWL<7293> A_IWL<7292> A_IWL<7291> A_IWL<7290> A_IWL<7289> A_IWL<7288> A_IWL<7287> A_IWL<7286> A_IWL<7285> A_IWL<7284> A_IWL<7283> A_IWL<7282> A_IWL<7281> A_IWL<7280> A_IWL<7279> A_IWL<7278> A_IWL<7277> A_IWL<7276> A_IWL<7275> A_IWL<7274> A_IWL<7273> A_IWL<7272> A_IWL<7271> A_IWL<7270> A_IWL<7269> A_IWL<7268> A_IWL<7267> A_IWL<7266> A_IWL<7265> A_IWL<7264> A_IWL<7263> A_IWL<7262> A_IWL<7261> A_IWL<7260> A_IWL<7259> A_IWL<7258> A_IWL<7257> A_IWL<7256> A_IWL<7255> A_IWL<7254> A_IWL<7253> A_IWL<7252> A_IWL<7251> A_IWL<7250> A_IWL<7249> A_IWL<7248> A_IWL<7247> A_IWL<7246> A_IWL<7245> A_IWL<7244> A_IWL<7243> A_IWL<7242> A_IWL<7241> A_IWL<7240> A_IWL<7239> A_IWL<7238> A_IWL<7237> A_IWL<7236> A_IWL<7235> A_IWL<7234> A_IWL<7233> A_IWL<7232> A_IWL<7231> A_IWL<7230> A_IWL<7229> A_IWL<7228> A_IWL<7227> A_IWL<7226> A_IWL<7225> A_IWL<7224> A_IWL<7223> A_IWL<7222> A_IWL<7221> A_IWL<7220> A_IWL<7219> A_IWL<7218> A_IWL<7217> A_IWL<7216> A_IWL<7215> A_IWL<7214> A_IWL<7213> A_IWL<7212> A_IWL<7211> A_IWL<7210> A_IWL<7209> A_IWL<7208> A_IWL<7207> A_IWL<7206> A_IWL<7205> A_IWL<7204> A_IWL<7203> A_IWL<7202> A_IWL<7201> A_IWL<7200> A_IWL<7199> A_IWL<7198> A_IWL<7197> A_IWL<7196> A_IWL<7195> A_IWL<7194> A_IWL<7193> A_IWL<7192> A_IWL<7191> A_IWL<7190> A_IWL<7189> A_IWL<7188> A_IWL<7187> A_IWL<7186> A_IWL<7185> A_IWL<7184> A_IWL<7183> A_IWL<7182> A_IWL<7181> A_IWL<7180> A_IWL<7179> A_IWL<7178> A_IWL<7177> A_IWL<7176> A_IWL<7175> A_IWL<7174> A_IWL<7173> A_IWL<7172> A_IWL<7171> A_IWL<7170> A_IWL<7169> A_IWL<7168> A_IWL<8191> A_IWL<8190> A_IWL<8189> A_IWL<8188> A_IWL<8187> A_IWL<8186> A_IWL<8185> A_IWL<8184> A_IWL<8183> A_IWL<8182> A_IWL<8181> A_IWL<8180> A_IWL<8179> A_IWL<8178> A_IWL<8177> A_IWL<8176> A_IWL<8175> A_IWL<8174> A_IWL<8173> A_IWL<8172> A_IWL<8171> A_IWL<8170> A_IWL<8169> A_IWL<8168> A_IWL<8167> A_IWL<8166> A_IWL<8165> A_IWL<8164> A_IWL<8163> A_IWL<8162> A_IWL<8161> A_IWL<8160> A_IWL<8159> A_IWL<8158> A_IWL<8157> A_IWL<8156> A_IWL<8155> A_IWL<8154> A_IWL<8153> A_IWL<8152> A_IWL<8151> A_IWL<8150> A_IWL<8149> A_IWL<8148> A_IWL<8147> A_IWL<8146> A_IWL<8145> A_IWL<8144> A_IWL<8143> A_IWL<8142> A_IWL<8141> A_IWL<8140> A_IWL<8139> A_IWL<8138> A_IWL<8137> A_IWL<8136> A_IWL<8135> A_IWL<8134> A_IWL<8133> A_IWL<8132> A_IWL<8131> A_IWL<8130> A_IWL<8129> A_IWL<8128> A_IWL<8127> A_IWL<8126> A_IWL<8125> A_IWL<8124> A_IWL<8123> A_IWL<8122> A_IWL<8121> A_IWL<8120> A_IWL<8119> A_IWL<8118> A_IWL<8117> A_IWL<8116> A_IWL<8115> A_IWL<8114> A_IWL<8113> A_IWL<8112> A_IWL<8111> A_IWL<8110> A_IWL<8109> A_IWL<8108> A_IWL<8107> A_IWL<8106> A_IWL<8105> A_IWL<8104> A_IWL<8103> A_IWL<8102> A_IWL<8101> A_IWL<8100> A_IWL<8099> A_IWL<8098> A_IWL<8097> A_IWL<8096> A_IWL<8095> A_IWL<8094> A_IWL<8093> A_IWL<8092> A_IWL<8091> A_IWL<8090> A_IWL<8089> A_IWL<8088> A_IWL<8087> A_IWL<8086> A_IWL<8085> A_IWL<8084> A_IWL<8083> A_IWL<8082> A_IWL<8081> A_IWL<8080> A_IWL<8079> A_IWL<8078> A_IWL<8077> A_IWL<8076> A_IWL<8075> A_IWL<8074> A_IWL<8073> A_IWL<8072> A_IWL<8071> A_IWL<8070> A_IWL<8069> A_IWL<8068> A_IWL<8067> A_IWL<8066> A_IWL<8065> A_IWL<8064> A_IWL<8063> A_IWL<8062> A_IWL<8061> A_IWL<8060> A_IWL<8059> A_IWL<8058> A_IWL<8057> A_IWL<8056> A_IWL<8055> A_IWL<8054> A_IWL<8053> A_IWL<8052> A_IWL<8051> A_IWL<8050> A_IWL<8049> A_IWL<8048> A_IWL<8047> A_IWL<8046> A_IWL<8045> A_IWL<8044> A_IWL<8043> A_IWL<8042> A_IWL<8041> A_IWL<8040> A_IWL<8039> A_IWL<8038> A_IWL<8037> A_IWL<8036> A_IWL<8035> A_IWL<8034> A_IWL<8033> A_IWL<8032> A_IWL<8031> A_IWL<8030> A_IWL<8029> A_IWL<8028> A_IWL<8027> A_IWL<8026> A_IWL<8025> A_IWL<8024> A_IWL<8023> A_IWL<8022> A_IWL<8021> A_IWL<8020> A_IWL<8019> A_IWL<8018> A_IWL<8017> A_IWL<8016> A_IWL<8015> A_IWL<8014> A_IWL<8013> A_IWL<8012> A_IWL<8011> A_IWL<8010> A_IWL<8009> A_IWL<8008> A_IWL<8007> A_IWL<8006> A_IWL<8005> A_IWL<8004> A_IWL<8003> A_IWL<8002> A_IWL<8001> A_IWL<8000> A_IWL<7999> A_IWL<7998> A_IWL<7997> A_IWL<7996> A_IWL<7995> A_IWL<7994> A_IWL<7993> A_IWL<7992> A_IWL<7991> A_IWL<7990> A_IWL<7989> A_IWL<7988> A_IWL<7987> A_IWL<7986> A_IWL<7985> A_IWL<7984> A_IWL<7983> A_IWL<7982> A_IWL<7981> A_IWL<7980> A_IWL<7979> A_IWL<7978> A_IWL<7977> A_IWL<7976> A_IWL<7975> A_IWL<7974> A_IWL<7973> A_IWL<7972> A_IWL<7971> A_IWL<7970> A_IWL<7969> A_IWL<7968> A_IWL<7967> A_IWL<7966> A_IWL<7965> A_IWL<7964> A_IWL<7963> A_IWL<7962> A_IWL<7961> A_IWL<7960> A_IWL<7959> A_IWL<7958> A_IWL<7957> A_IWL<7956> A_IWL<7955> A_IWL<7954> A_IWL<7953> A_IWL<7952> A_IWL<7951> A_IWL<7950> A_IWL<7949> A_IWL<7948> A_IWL<7947> A_IWL<7946> A_IWL<7945> A_IWL<7944> A_IWL<7943> A_IWL<7942> A_IWL<7941> A_IWL<7940> A_IWL<7939> A_IWL<7938> A_IWL<7937> A_IWL<7936> A_IWL<7935> A_IWL<7934> A_IWL<7933> A_IWL<7932> A_IWL<7931> A_IWL<7930> A_IWL<7929> A_IWL<7928> A_IWL<7927> A_IWL<7926> A_IWL<7925> A_IWL<7924> A_IWL<7923> A_IWL<7922> A_IWL<7921> A_IWL<7920> A_IWL<7919> A_IWL<7918> A_IWL<7917> A_IWL<7916> A_IWL<7915> A_IWL<7914> A_IWL<7913> A_IWL<7912> A_IWL<7911> A_IWL<7910> A_IWL<7909> A_IWL<7908> A_IWL<7907> A_IWL<7906> A_IWL<7905> A_IWL<7904> A_IWL<7903> A_IWL<7902> A_IWL<7901> A_IWL<7900> A_IWL<7899> A_IWL<7898> A_IWL<7897> A_IWL<7896> A_IWL<7895> A_IWL<7894> A_IWL<7893> A_IWL<7892> A_IWL<7891> A_IWL<7890> A_IWL<7889> A_IWL<7888> A_IWL<7887> A_IWL<7886> A_IWL<7885> A_IWL<7884> A_IWL<7883> A_IWL<7882> A_IWL<7881> A_IWL<7880> A_IWL<7879> A_IWL<7878> A_IWL<7877> A_IWL<7876> A_IWL<7875> A_IWL<7874> A_IWL<7873> A_IWL<7872> A_IWL<7871> A_IWL<7870> A_IWL<7869> A_IWL<7868> A_IWL<7867> A_IWL<7866> A_IWL<7865> A_IWL<7864> A_IWL<7863> A_IWL<7862> A_IWL<7861> A_IWL<7860> A_IWL<7859> A_IWL<7858> A_IWL<7857> A_IWL<7856> A_IWL<7855> A_IWL<7854> A_IWL<7853> A_IWL<7852> A_IWL<7851> A_IWL<7850> A_IWL<7849> A_IWL<7848> A_IWL<7847> A_IWL<7846> A_IWL<7845> A_IWL<7844> A_IWL<7843> A_IWL<7842> A_IWL<7841> A_IWL<7840> A_IWL<7839> A_IWL<7838> A_IWL<7837> A_IWL<7836> A_IWL<7835> A_IWL<7834> A_IWL<7833> A_IWL<7832> A_IWL<7831> A_IWL<7830> A_IWL<7829> A_IWL<7828> A_IWL<7827> A_IWL<7826> A_IWL<7825> A_IWL<7824> A_IWL<7823> A_IWL<7822> A_IWL<7821> A_IWL<7820> A_IWL<7819> A_IWL<7818> A_IWL<7817> A_IWL<7816> A_IWL<7815> A_IWL<7814> A_IWL<7813> A_IWL<7812> A_IWL<7811> A_IWL<7810> A_IWL<7809> A_IWL<7808> A_IWL<7807> A_IWL<7806> A_IWL<7805> A_IWL<7804> A_IWL<7803> A_IWL<7802> A_IWL<7801> A_IWL<7800> A_IWL<7799> A_IWL<7798> A_IWL<7797> A_IWL<7796> A_IWL<7795> A_IWL<7794> A_IWL<7793> A_IWL<7792> A_IWL<7791> A_IWL<7790> A_IWL<7789> A_IWL<7788> A_IWL<7787> A_IWL<7786> A_IWL<7785> A_IWL<7784> A_IWL<7783> A_IWL<7782> A_IWL<7781> A_IWL<7780> A_IWL<7779> A_IWL<7778> A_IWL<7777> A_IWL<7776> A_IWL<7775> A_IWL<7774> A_IWL<7773> A_IWL<7772> A_IWL<7771> A_IWL<7770> A_IWL<7769> A_IWL<7768> A_IWL<7767> A_IWL<7766> A_IWL<7765> A_IWL<7764> A_IWL<7763> A_IWL<7762> A_IWL<7761> A_IWL<7760> A_IWL<7759> A_IWL<7758> A_IWL<7757> A_IWL<7756> A_IWL<7755> A_IWL<7754> A_IWL<7753> A_IWL<7752> A_IWL<7751> A_IWL<7750> A_IWL<7749> A_IWL<7748> A_IWL<7747> A_IWL<7746> A_IWL<7745> A_IWL<7744> A_IWL<7743> A_IWL<7742> A_IWL<7741> A_IWL<7740> A_IWL<7739> A_IWL<7738> A_IWL<7737> A_IWL<7736> A_IWL<7735> A_IWL<7734> A_IWL<7733> A_IWL<7732> A_IWL<7731> A_IWL<7730> A_IWL<7729> A_IWL<7728> A_IWL<7727> A_IWL<7726> A_IWL<7725> A_IWL<7724> A_IWL<7723> A_IWL<7722> A_IWL<7721> A_IWL<7720> A_IWL<7719> A_IWL<7718> A_IWL<7717> A_IWL<7716> A_IWL<7715> A_IWL<7714> A_IWL<7713> A_IWL<7712> A_IWL<7711> A_IWL<7710> A_IWL<7709> A_IWL<7708> A_IWL<7707> A_IWL<7706> A_IWL<7705> A_IWL<7704> A_IWL<7703> A_IWL<7702> A_IWL<7701> A_IWL<7700> A_IWL<7699> A_IWL<7698> A_IWL<7697> A_IWL<7696> A_IWL<7695> A_IWL<7694> A_IWL<7693> A_IWL<7692> A_IWL<7691> A_IWL<7690> A_IWL<7689> A_IWL<7688> A_IWL<7687> A_IWL<7686> A_IWL<7685> A_IWL<7684> A_IWL<7683> A_IWL<7682> A_IWL<7681> A_IWL<7680> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<14> A_BLC<29> A_BLC<28> A_BLC_TOP<29> A_BLC_TOP<28> A_BLT<29> A_BLT<28> A_BLT_TOP<29> A_BLT_TOP<28> A_IWL<7167> A_IWL<7166> A_IWL<7165> A_IWL<7164> A_IWL<7163> A_IWL<7162> A_IWL<7161> A_IWL<7160> A_IWL<7159> A_IWL<7158> A_IWL<7157> A_IWL<7156> A_IWL<7155> A_IWL<7154> A_IWL<7153> A_IWL<7152> A_IWL<7151> A_IWL<7150> A_IWL<7149> A_IWL<7148> A_IWL<7147> A_IWL<7146> A_IWL<7145> A_IWL<7144> A_IWL<7143> A_IWL<7142> A_IWL<7141> A_IWL<7140> A_IWL<7139> A_IWL<7138> A_IWL<7137> A_IWL<7136> A_IWL<7135> A_IWL<7134> A_IWL<7133> A_IWL<7132> A_IWL<7131> A_IWL<7130> A_IWL<7129> A_IWL<7128> A_IWL<7127> A_IWL<7126> A_IWL<7125> A_IWL<7124> A_IWL<7123> A_IWL<7122> A_IWL<7121> A_IWL<7120> A_IWL<7119> A_IWL<7118> A_IWL<7117> A_IWL<7116> A_IWL<7115> A_IWL<7114> A_IWL<7113> A_IWL<7112> A_IWL<7111> A_IWL<7110> A_IWL<7109> A_IWL<7108> A_IWL<7107> A_IWL<7106> A_IWL<7105> A_IWL<7104> A_IWL<7103> A_IWL<7102> A_IWL<7101> A_IWL<7100> A_IWL<7099> A_IWL<7098> A_IWL<7097> A_IWL<7096> A_IWL<7095> A_IWL<7094> A_IWL<7093> A_IWL<7092> A_IWL<7091> A_IWL<7090> A_IWL<7089> A_IWL<7088> A_IWL<7087> A_IWL<7086> A_IWL<7085> A_IWL<7084> A_IWL<7083> A_IWL<7082> A_IWL<7081> A_IWL<7080> A_IWL<7079> A_IWL<7078> A_IWL<7077> A_IWL<7076> A_IWL<7075> A_IWL<7074> A_IWL<7073> A_IWL<7072> A_IWL<7071> A_IWL<7070> A_IWL<7069> A_IWL<7068> A_IWL<7067> A_IWL<7066> A_IWL<7065> A_IWL<7064> A_IWL<7063> A_IWL<7062> A_IWL<7061> A_IWL<7060> A_IWL<7059> A_IWL<7058> A_IWL<7057> A_IWL<7056> A_IWL<7055> A_IWL<7054> A_IWL<7053> A_IWL<7052> A_IWL<7051> A_IWL<7050> A_IWL<7049> A_IWL<7048> A_IWL<7047> A_IWL<7046> A_IWL<7045> A_IWL<7044> A_IWL<7043> A_IWL<7042> A_IWL<7041> A_IWL<7040> A_IWL<7039> A_IWL<7038> A_IWL<7037> A_IWL<7036> A_IWL<7035> A_IWL<7034> A_IWL<7033> A_IWL<7032> A_IWL<7031> A_IWL<7030> A_IWL<7029> A_IWL<7028> A_IWL<7027> A_IWL<7026> A_IWL<7025> A_IWL<7024> A_IWL<7023> A_IWL<7022> A_IWL<7021> A_IWL<7020> A_IWL<7019> A_IWL<7018> A_IWL<7017> A_IWL<7016> A_IWL<7015> A_IWL<7014> A_IWL<7013> A_IWL<7012> A_IWL<7011> A_IWL<7010> A_IWL<7009> A_IWL<7008> A_IWL<7007> A_IWL<7006> A_IWL<7005> A_IWL<7004> A_IWL<7003> A_IWL<7002> A_IWL<7001> A_IWL<7000> A_IWL<6999> A_IWL<6998> A_IWL<6997> A_IWL<6996> A_IWL<6995> A_IWL<6994> A_IWL<6993> A_IWL<6992> A_IWL<6991> A_IWL<6990> A_IWL<6989> A_IWL<6988> A_IWL<6987> A_IWL<6986> A_IWL<6985> A_IWL<6984> A_IWL<6983> A_IWL<6982> A_IWL<6981> A_IWL<6980> A_IWL<6979> A_IWL<6978> A_IWL<6977> A_IWL<6976> A_IWL<6975> A_IWL<6974> A_IWL<6973> A_IWL<6972> A_IWL<6971> A_IWL<6970> A_IWL<6969> A_IWL<6968> A_IWL<6967> A_IWL<6966> A_IWL<6965> A_IWL<6964> A_IWL<6963> A_IWL<6962> A_IWL<6961> A_IWL<6960> A_IWL<6959> A_IWL<6958> A_IWL<6957> A_IWL<6956> A_IWL<6955> A_IWL<6954> A_IWL<6953> A_IWL<6952> A_IWL<6951> A_IWL<6950> A_IWL<6949> A_IWL<6948> A_IWL<6947> A_IWL<6946> A_IWL<6945> A_IWL<6944> A_IWL<6943> A_IWL<6942> A_IWL<6941> A_IWL<6940> A_IWL<6939> A_IWL<6938> A_IWL<6937> A_IWL<6936> A_IWL<6935> A_IWL<6934> A_IWL<6933> A_IWL<6932> A_IWL<6931> A_IWL<6930> A_IWL<6929> A_IWL<6928> A_IWL<6927> A_IWL<6926> A_IWL<6925> A_IWL<6924> A_IWL<6923> A_IWL<6922> A_IWL<6921> A_IWL<6920> A_IWL<6919> A_IWL<6918> A_IWL<6917> A_IWL<6916> A_IWL<6915> A_IWL<6914> A_IWL<6913> A_IWL<6912> A_IWL<6911> A_IWL<6910> A_IWL<6909> A_IWL<6908> A_IWL<6907> A_IWL<6906> A_IWL<6905> A_IWL<6904> A_IWL<6903> A_IWL<6902> A_IWL<6901> A_IWL<6900> A_IWL<6899> A_IWL<6898> A_IWL<6897> A_IWL<6896> A_IWL<6895> A_IWL<6894> A_IWL<6893> A_IWL<6892> A_IWL<6891> A_IWL<6890> A_IWL<6889> A_IWL<6888> A_IWL<6887> A_IWL<6886> A_IWL<6885> A_IWL<6884> A_IWL<6883> A_IWL<6882> A_IWL<6881> A_IWL<6880> A_IWL<6879> A_IWL<6878> A_IWL<6877> A_IWL<6876> A_IWL<6875> A_IWL<6874> A_IWL<6873> A_IWL<6872> A_IWL<6871> A_IWL<6870> A_IWL<6869> A_IWL<6868> A_IWL<6867> A_IWL<6866> A_IWL<6865> A_IWL<6864> A_IWL<6863> A_IWL<6862> A_IWL<6861> A_IWL<6860> A_IWL<6859> A_IWL<6858> A_IWL<6857> A_IWL<6856> A_IWL<6855> A_IWL<6854> A_IWL<6853> A_IWL<6852> A_IWL<6851> A_IWL<6850> A_IWL<6849> A_IWL<6848> A_IWL<6847> A_IWL<6846> A_IWL<6845> A_IWL<6844> A_IWL<6843> A_IWL<6842> A_IWL<6841> A_IWL<6840> A_IWL<6839> A_IWL<6838> A_IWL<6837> A_IWL<6836> A_IWL<6835> A_IWL<6834> A_IWL<6833> A_IWL<6832> A_IWL<6831> A_IWL<6830> A_IWL<6829> A_IWL<6828> A_IWL<6827> A_IWL<6826> A_IWL<6825> A_IWL<6824> A_IWL<6823> A_IWL<6822> A_IWL<6821> A_IWL<6820> A_IWL<6819> A_IWL<6818> A_IWL<6817> A_IWL<6816> A_IWL<6815> A_IWL<6814> A_IWL<6813> A_IWL<6812> A_IWL<6811> A_IWL<6810> A_IWL<6809> A_IWL<6808> A_IWL<6807> A_IWL<6806> A_IWL<6805> A_IWL<6804> A_IWL<6803> A_IWL<6802> A_IWL<6801> A_IWL<6800> A_IWL<6799> A_IWL<6798> A_IWL<6797> A_IWL<6796> A_IWL<6795> A_IWL<6794> A_IWL<6793> A_IWL<6792> A_IWL<6791> A_IWL<6790> A_IWL<6789> A_IWL<6788> A_IWL<6787> A_IWL<6786> A_IWL<6785> A_IWL<6784> A_IWL<6783> A_IWL<6782> A_IWL<6781> A_IWL<6780> A_IWL<6779> A_IWL<6778> A_IWL<6777> A_IWL<6776> A_IWL<6775> A_IWL<6774> A_IWL<6773> A_IWL<6772> A_IWL<6771> A_IWL<6770> A_IWL<6769> A_IWL<6768> A_IWL<6767> A_IWL<6766> A_IWL<6765> A_IWL<6764> A_IWL<6763> A_IWL<6762> A_IWL<6761> A_IWL<6760> A_IWL<6759> A_IWL<6758> A_IWL<6757> A_IWL<6756> A_IWL<6755> A_IWL<6754> A_IWL<6753> A_IWL<6752> A_IWL<6751> A_IWL<6750> A_IWL<6749> A_IWL<6748> A_IWL<6747> A_IWL<6746> A_IWL<6745> A_IWL<6744> A_IWL<6743> A_IWL<6742> A_IWL<6741> A_IWL<6740> A_IWL<6739> A_IWL<6738> A_IWL<6737> A_IWL<6736> A_IWL<6735> A_IWL<6734> A_IWL<6733> A_IWL<6732> A_IWL<6731> A_IWL<6730> A_IWL<6729> A_IWL<6728> A_IWL<6727> A_IWL<6726> A_IWL<6725> A_IWL<6724> A_IWL<6723> A_IWL<6722> A_IWL<6721> A_IWL<6720> A_IWL<6719> A_IWL<6718> A_IWL<6717> A_IWL<6716> A_IWL<6715> A_IWL<6714> A_IWL<6713> A_IWL<6712> A_IWL<6711> A_IWL<6710> A_IWL<6709> A_IWL<6708> A_IWL<6707> A_IWL<6706> A_IWL<6705> A_IWL<6704> A_IWL<6703> A_IWL<6702> A_IWL<6701> A_IWL<6700> A_IWL<6699> A_IWL<6698> A_IWL<6697> A_IWL<6696> A_IWL<6695> A_IWL<6694> A_IWL<6693> A_IWL<6692> A_IWL<6691> A_IWL<6690> A_IWL<6689> A_IWL<6688> A_IWL<6687> A_IWL<6686> A_IWL<6685> A_IWL<6684> A_IWL<6683> A_IWL<6682> A_IWL<6681> A_IWL<6680> A_IWL<6679> A_IWL<6678> A_IWL<6677> A_IWL<6676> A_IWL<6675> A_IWL<6674> A_IWL<6673> A_IWL<6672> A_IWL<6671> A_IWL<6670> A_IWL<6669> A_IWL<6668> A_IWL<6667> A_IWL<6666> A_IWL<6665> A_IWL<6664> A_IWL<6663> A_IWL<6662> A_IWL<6661> A_IWL<6660> A_IWL<6659> A_IWL<6658> A_IWL<6657> A_IWL<6656> A_IWL<7679> A_IWL<7678> A_IWL<7677> A_IWL<7676> A_IWL<7675> A_IWL<7674> A_IWL<7673> A_IWL<7672> A_IWL<7671> A_IWL<7670> A_IWL<7669> A_IWL<7668> A_IWL<7667> A_IWL<7666> A_IWL<7665> A_IWL<7664> A_IWL<7663> A_IWL<7662> A_IWL<7661> A_IWL<7660> A_IWL<7659> A_IWL<7658> A_IWL<7657> A_IWL<7656> A_IWL<7655> A_IWL<7654> A_IWL<7653> A_IWL<7652> A_IWL<7651> A_IWL<7650> A_IWL<7649> A_IWL<7648> A_IWL<7647> A_IWL<7646> A_IWL<7645> A_IWL<7644> A_IWL<7643> A_IWL<7642> A_IWL<7641> A_IWL<7640> A_IWL<7639> A_IWL<7638> A_IWL<7637> A_IWL<7636> A_IWL<7635> A_IWL<7634> A_IWL<7633> A_IWL<7632> A_IWL<7631> A_IWL<7630> A_IWL<7629> A_IWL<7628> A_IWL<7627> A_IWL<7626> A_IWL<7625> A_IWL<7624> A_IWL<7623> A_IWL<7622> A_IWL<7621> A_IWL<7620> A_IWL<7619> A_IWL<7618> A_IWL<7617> A_IWL<7616> A_IWL<7615> A_IWL<7614> A_IWL<7613> A_IWL<7612> A_IWL<7611> A_IWL<7610> A_IWL<7609> A_IWL<7608> A_IWL<7607> A_IWL<7606> A_IWL<7605> A_IWL<7604> A_IWL<7603> A_IWL<7602> A_IWL<7601> A_IWL<7600> A_IWL<7599> A_IWL<7598> A_IWL<7597> A_IWL<7596> A_IWL<7595> A_IWL<7594> A_IWL<7593> A_IWL<7592> A_IWL<7591> A_IWL<7590> A_IWL<7589> A_IWL<7588> A_IWL<7587> A_IWL<7586> A_IWL<7585> A_IWL<7584> A_IWL<7583> A_IWL<7582> A_IWL<7581> A_IWL<7580> A_IWL<7579> A_IWL<7578> A_IWL<7577> A_IWL<7576> A_IWL<7575> A_IWL<7574> A_IWL<7573> A_IWL<7572> A_IWL<7571> A_IWL<7570> A_IWL<7569> A_IWL<7568> A_IWL<7567> A_IWL<7566> A_IWL<7565> A_IWL<7564> A_IWL<7563> A_IWL<7562> A_IWL<7561> A_IWL<7560> A_IWL<7559> A_IWL<7558> A_IWL<7557> A_IWL<7556> A_IWL<7555> A_IWL<7554> A_IWL<7553> A_IWL<7552> A_IWL<7551> A_IWL<7550> A_IWL<7549> A_IWL<7548> A_IWL<7547> A_IWL<7546> A_IWL<7545> A_IWL<7544> A_IWL<7543> A_IWL<7542> A_IWL<7541> A_IWL<7540> A_IWL<7539> A_IWL<7538> A_IWL<7537> A_IWL<7536> A_IWL<7535> A_IWL<7534> A_IWL<7533> A_IWL<7532> A_IWL<7531> A_IWL<7530> A_IWL<7529> A_IWL<7528> A_IWL<7527> A_IWL<7526> A_IWL<7525> A_IWL<7524> A_IWL<7523> A_IWL<7522> A_IWL<7521> A_IWL<7520> A_IWL<7519> A_IWL<7518> A_IWL<7517> A_IWL<7516> A_IWL<7515> A_IWL<7514> A_IWL<7513> A_IWL<7512> A_IWL<7511> A_IWL<7510> A_IWL<7509> A_IWL<7508> A_IWL<7507> A_IWL<7506> A_IWL<7505> A_IWL<7504> A_IWL<7503> A_IWL<7502> A_IWL<7501> A_IWL<7500> A_IWL<7499> A_IWL<7498> A_IWL<7497> A_IWL<7496> A_IWL<7495> A_IWL<7494> A_IWL<7493> A_IWL<7492> A_IWL<7491> A_IWL<7490> A_IWL<7489> A_IWL<7488> A_IWL<7487> A_IWL<7486> A_IWL<7485> A_IWL<7484> A_IWL<7483> A_IWL<7482> A_IWL<7481> A_IWL<7480> A_IWL<7479> A_IWL<7478> A_IWL<7477> A_IWL<7476> A_IWL<7475> A_IWL<7474> A_IWL<7473> A_IWL<7472> A_IWL<7471> A_IWL<7470> A_IWL<7469> A_IWL<7468> A_IWL<7467> A_IWL<7466> A_IWL<7465> A_IWL<7464> A_IWL<7463> A_IWL<7462> A_IWL<7461> A_IWL<7460> A_IWL<7459> A_IWL<7458> A_IWL<7457> A_IWL<7456> A_IWL<7455> A_IWL<7454> A_IWL<7453> A_IWL<7452> A_IWL<7451> A_IWL<7450> A_IWL<7449> A_IWL<7448> A_IWL<7447> A_IWL<7446> A_IWL<7445> A_IWL<7444> A_IWL<7443> A_IWL<7442> A_IWL<7441> A_IWL<7440> A_IWL<7439> A_IWL<7438> A_IWL<7437> A_IWL<7436> A_IWL<7435> A_IWL<7434> A_IWL<7433> A_IWL<7432> A_IWL<7431> A_IWL<7430> A_IWL<7429> A_IWL<7428> A_IWL<7427> A_IWL<7426> A_IWL<7425> A_IWL<7424> A_IWL<7423> A_IWL<7422> A_IWL<7421> A_IWL<7420> A_IWL<7419> A_IWL<7418> A_IWL<7417> A_IWL<7416> A_IWL<7415> A_IWL<7414> A_IWL<7413> A_IWL<7412> A_IWL<7411> A_IWL<7410> A_IWL<7409> A_IWL<7408> A_IWL<7407> A_IWL<7406> A_IWL<7405> A_IWL<7404> A_IWL<7403> A_IWL<7402> A_IWL<7401> A_IWL<7400> A_IWL<7399> A_IWL<7398> A_IWL<7397> A_IWL<7396> A_IWL<7395> A_IWL<7394> A_IWL<7393> A_IWL<7392> A_IWL<7391> A_IWL<7390> A_IWL<7389> A_IWL<7388> A_IWL<7387> A_IWL<7386> A_IWL<7385> A_IWL<7384> A_IWL<7383> A_IWL<7382> A_IWL<7381> A_IWL<7380> A_IWL<7379> A_IWL<7378> A_IWL<7377> A_IWL<7376> A_IWL<7375> A_IWL<7374> A_IWL<7373> A_IWL<7372> A_IWL<7371> A_IWL<7370> A_IWL<7369> A_IWL<7368> A_IWL<7367> A_IWL<7366> A_IWL<7365> A_IWL<7364> A_IWL<7363> A_IWL<7362> A_IWL<7361> A_IWL<7360> A_IWL<7359> A_IWL<7358> A_IWL<7357> A_IWL<7356> A_IWL<7355> A_IWL<7354> A_IWL<7353> A_IWL<7352> A_IWL<7351> A_IWL<7350> A_IWL<7349> A_IWL<7348> A_IWL<7347> A_IWL<7346> A_IWL<7345> A_IWL<7344> A_IWL<7343> A_IWL<7342> A_IWL<7341> A_IWL<7340> A_IWL<7339> A_IWL<7338> A_IWL<7337> A_IWL<7336> A_IWL<7335> A_IWL<7334> A_IWL<7333> A_IWL<7332> A_IWL<7331> A_IWL<7330> A_IWL<7329> A_IWL<7328> A_IWL<7327> A_IWL<7326> A_IWL<7325> A_IWL<7324> A_IWL<7323> A_IWL<7322> A_IWL<7321> A_IWL<7320> A_IWL<7319> A_IWL<7318> A_IWL<7317> A_IWL<7316> A_IWL<7315> A_IWL<7314> A_IWL<7313> A_IWL<7312> A_IWL<7311> A_IWL<7310> A_IWL<7309> A_IWL<7308> A_IWL<7307> A_IWL<7306> A_IWL<7305> A_IWL<7304> A_IWL<7303> A_IWL<7302> A_IWL<7301> A_IWL<7300> A_IWL<7299> A_IWL<7298> A_IWL<7297> A_IWL<7296> A_IWL<7295> A_IWL<7294> A_IWL<7293> A_IWL<7292> A_IWL<7291> A_IWL<7290> A_IWL<7289> A_IWL<7288> A_IWL<7287> A_IWL<7286> A_IWL<7285> A_IWL<7284> A_IWL<7283> A_IWL<7282> A_IWL<7281> A_IWL<7280> A_IWL<7279> A_IWL<7278> A_IWL<7277> A_IWL<7276> A_IWL<7275> A_IWL<7274> A_IWL<7273> A_IWL<7272> A_IWL<7271> A_IWL<7270> A_IWL<7269> A_IWL<7268> A_IWL<7267> A_IWL<7266> A_IWL<7265> A_IWL<7264> A_IWL<7263> A_IWL<7262> A_IWL<7261> A_IWL<7260> A_IWL<7259> A_IWL<7258> A_IWL<7257> A_IWL<7256> A_IWL<7255> A_IWL<7254> A_IWL<7253> A_IWL<7252> A_IWL<7251> A_IWL<7250> A_IWL<7249> A_IWL<7248> A_IWL<7247> A_IWL<7246> A_IWL<7245> A_IWL<7244> A_IWL<7243> A_IWL<7242> A_IWL<7241> A_IWL<7240> A_IWL<7239> A_IWL<7238> A_IWL<7237> A_IWL<7236> A_IWL<7235> A_IWL<7234> A_IWL<7233> A_IWL<7232> A_IWL<7231> A_IWL<7230> A_IWL<7229> A_IWL<7228> A_IWL<7227> A_IWL<7226> A_IWL<7225> A_IWL<7224> A_IWL<7223> A_IWL<7222> A_IWL<7221> A_IWL<7220> A_IWL<7219> A_IWL<7218> A_IWL<7217> A_IWL<7216> A_IWL<7215> A_IWL<7214> A_IWL<7213> A_IWL<7212> A_IWL<7211> A_IWL<7210> A_IWL<7209> A_IWL<7208> A_IWL<7207> A_IWL<7206> A_IWL<7205> A_IWL<7204> A_IWL<7203> A_IWL<7202> A_IWL<7201> A_IWL<7200> A_IWL<7199> A_IWL<7198> A_IWL<7197> A_IWL<7196> A_IWL<7195> A_IWL<7194> A_IWL<7193> A_IWL<7192> A_IWL<7191> A_IWL<7190> A_IWL<7189> A_IWL<7188> A_IWL<7187> A_IWL<7186> A_IWL<7185> A_IWL<7184> A_IWL<7183> A_IWL<7182> A_IWL<7181> A_IWL<7180> A_IWL<7179> A_IWL<7178> A_IWL<7177> A_IWL<7176> A_IWL<7175> A_IWL<7174> A_IWL<7173> A_IWL<7172> A_IWL<7171> A_IWL<7170> A_IWL<7169> A_IWL<7168> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<13> A_BLC<27> A_BLC<26> A_BLC_TOP<27> A_BLC_TOP<26> A_BLT<27> A_BLT<26> A_BLT_TOP<27> A_BLT_TOP<26> A_IWL<6655> A_IWL<6654> A_IWL<6653> A_IWL<6652> A_IWL<6651> A_IWL<6650> A_IWL<6649> A_IWL<6648> A_IWL<6647> A_IWL<6646> A_IWL<6645> A_IWL<6644> A_IWL<6643> A_IWL<6642> A_IWL<6641> A_IWL<6640> A_IWL<6639> A_IWL<6638> A_IWL<6637> A_IWL<6636> A_IWL<6635> A_IWL<6634> A_IWL<6633> A_IWL<6632> A_IWL<6631> A_IWL<6630> A_IWL<6629> A_IWL<6628> A_IWL<6627> A_IWL<6626> A_IWL<6625> A_IWL<6624> A_IWL<6623> A_IWL<6622> A_IWL<6621> A_IWL<6620> A_IWL<6619> A_IWL<6618> A_IWL<6617> A_IWL<6616> A_IWL<6615> A_IWL<6614> A_IWL<6613> A_IWL<6612> A_IWL<6611> A_IWL<6610> A_IWL<6609> A_IWL<6608> A_IWL<6607> A_IWL<6606> A_IWL<6605> A_IWL<6604> A_IWL<6603> A_IWL<6602> A_IWL<6601> A_IWL<6600> A_IWL<6599> A_IWL<6598> A_IWL<6597> A_IWL<6596> A_IWL<6595> A_IWL<6594> A_IWL<6593> A_IWL<6592> A_IWL<6591> A_IWL<6590> A_IWL<6589> A_IWL<6588> A_IWL<6587> A_IWL<6586> A_IWL<6585> A_IWL<6584> A_IWL<6583> A_IWL<6582> A_IWL<6581> A_IWL<6580> A_IWL<6579> A_IWL<6578> A_IWL<6577> A_IWL<6576> A_IWL<6575> A_IWL<6574> A_IWL<6573> A_IWL<6572> A_IWL<6571> A_IWL<6570> A_IWL<6569> A_IWL<6568> A_IWL<6567> A_IWL<6566> A_IWL<6565> A_IWL<6564> A_IWL<6563> A_IWL<6562> A_IWL<6561> A_IWL<6560> A_IWL<6559> A_IWL<6558> A_IWL<6557> A_IWL<6556> A_IWL<6555> A_IWL<6554> A_IWL<6553> A_IWL<6552> A_IWL<6551> A_IWL<6550> A_IWL<6549> A_IWL<6548> A_IWL<6547> A_IWL<6546> A_IWL<6545> A_IWL<6544> A_IWL<6543> A_IWL<6542> A_IWL<6541> A_IWL<6540> A_IWL<6539> A_IWL<6538> A_IWL<6537> A_IWL<6536> A_IWL<6535> A_IWL<6534> A_IWL<6533> A_IWL<6532> A_IWL<6531> A_IWL<6530> A_IWL<6529> A_IWL<6528> A_IWL<6527> A_IWL<6526> A_IWL<6525> A_IWL<6524> A_IWL<6523> A_IWL<6522> A_IWL<6521> A_IWL<6520> A_IWL<6519> A_IWL<6518> A_IWL<6517> A_IWL<6516> A_IWL<6515> A_IWL<6514> A_IWL<6513> A_IWL<6512> A_IWL<6511> A_IWL<6510> A_IWL<6509> A_IWL<6508> A_IWL<6507> A_IWL<6506> A_IWL<6505> A_IWL<6504> A_IWL<6503> A_IWL<6502> A_IWL<6501> A_IWL<6500> A_IWL<6499> A_IWL<6498> A_IWL<6497> A_IWL<6496> A_IWL<6495> A_IWL<6494> A_IWL<6493> A_IWL<6492> A_IWL<6491> A_IWL<6490> A_IWL<6489> A_IWL<6488> A_IWL<6487> A_IWL<6486> A_IWL<6485> A_IWL<6484> A_IWL<6483> A_IWL<6482> A_IWL<6481> A_IWL<6480> A_IWL<6479> A_IWL<6478> A_IWL<6477> A_IWL<6476> A_IWL<6475> A_IWL<6474> A_IWL<6473> A_IWL<6472> A_IWL<6471> A_IWL<6470> A_IWL<6469> A_IWL<6468> A_IWL<6467> A_IWL<6466> A_IWL<6465> A_IWL<6464> A_IWL<6463> A_IWL<6462> A_IWL<6461> A_IWL<6460> A_IWL<6459> A_IWL<6458> A_IWL<6457> A_IWL<6456> A_IWL<6455> A_IWL<6454> A_IWL<6453> A_IWL<6452> A_IWL<6451> A_IWL<6450> A_IWL<6449> A_IWL<6448> A_IWL<6447> A_IWL<6446> A_IWL<6445> A_IWL<6444> A_IWL<6443> A_IWL<6442> A_IWL<6441> A_IWL<6440> A_IWL<6439> A_IWL<6438> A_IWL<6437> A_IWL<6436> A_IWL<6435> A_IWL<6434> A_IWL<6433> A_IWL<6432> A_IWL<6431> A_IWL<6430> A_IWL<6429> A_IWL<6428> A_IWL<6427> A_IWL<6426> A_IWL<6425> A_IWL<6424> A_IWL<6423> A_IWL<6422> A_IWL<6421> A_IWL<6420> A_IWL<6419> A_IWL<6418> A_IWL<6417> A_IWL<6416> A_IWL<6415> A_IWL<6414> A_IWL<6413> A_IWL<6412> A_IWL<6411> A_IWL<6410> A_IWL<6409> A_IWL<6408> A_IWL<6407> A_IWL<6406> A_IWL<6405> A_IWL<6404> A_IWL<6403> A_IWL<6402> A_IWL<6401> A_IWL<6400> A_IWL<6399> A_IWL<6398> A_IWL<6397> A_IWL<6396> A_IWL<6395> A_IWL<6394> A_IWL<6393> A_IWL<6392> A_IWL<6391> A_IWL<6390> A_IWL<6389> A_IWL<6388> A_IWL<6387> A_IWL<6386> A_IWL<6385> A_IWL<6384> A_IWL<6383> A_IWL<6382> A_IWL<6381> A_IWL<6380> A_IWL<6379> A_IWL<6378> A_IWL<6377> A_IWL<6376> A_IWL<6375> A_IWL<6374> A_IWL<6373> A_IWL<6372> A_IWL<6371> A_IWL<6370> A_IWL<6369> A_IWL<6368> A_IWL<6367> A_IWL<6366> A_IWL<6365> A_IWL<6364> A_IWL<6363> A_IWL<6362> A_IWL<6361> A_IWL<6360> A_IWL<6359> A_IWL<6358> A_IWL<6357> A_IWL<6356> A_IWL<6355> A_IWL<6354> A_IWL<6353> A_IWL<6352> A_IWL<6351> A_IWL<6350> A_IWL<6349> A_IWL<6348> A_IWL<6347> A_IWL<6346> A_IWL<6345> A_IWL<6344> A_IWL<6343> A_IWL<6342> A_IWL<6341> A_IWL<6340> A_IWL<6339> A_IWL<6338> A_IWL<6337> A_IWL<6336> A_IWL<6335> A_IWL<6334> A_IWL<6333> A_IWL<6332> A_IWL<6331> A_IWL<6330> A_IWL<6329> A_IWL<6328> A_IWL<6327> A_IWL<6326> A_IWL<6325> A_IWL<6324> A_IWL<6323> A_IWL<6322> A_IWL<6321> A_IWL<6320> A_IWL<6319> A_IWL<6318> A_IWL<6317> A_IWL<6316> A_IWL<6315> A_IWL<6314> A_IWL<6313> A_IWL<6312> A_IWL<6311> A_IWL<6310> A_IWL<6309> A_IWL<6308> A_IWL<6307> A_IWL<6306> A_IWL<6305> A_IWL<6304> A_IWL<6303> A_IWL<6302> A_IWL<6301> A_IWL<6300> A_IWL<6299> A_IWL<6298> A_IWL<6297> A_IWL<6296> A_IWL<6295> A_IWL<6294> A_IWL<6293> A_IWL<6292> A_IWL<6291> A_IWL<6290> A_IWL<6289> A_IWL<6288> A_IWL<6287> A_IWL<6286> A_IWL<6285> A_IWL<6284> A_IWL<6283> A_IWL<6282> A_IWL<6281> A_IWL<6280> A_IWL<6279> A_IWL<6278> A_IWL<6277> A_IWL<6276> A_IWL<6275> A_IWL<6274> A_IWL<6273> A_IWL<6272> A_IWL<6271> A_IWL<6270> A_IWL<6269> A_IWL<6268> A_IWL<6267> A_IWL<6266> A_IWL<6265> A_IWL<6264> A_IWL<6263> A_IWL<6262> A_IWL<6261> A_IWL<6260> A_IWL<6259> A_IWL<6258> A_IWL<6257> A_IWL<6256> A_IWL<6255> A_IWL<6254> A_IWL<6253> A_IWL<6252> A_IWL<6251> A_IWL<6250> A_IWL<6249> A_IWL<6248> A_IWL<6247> A_IWL<6246> A_IWL<6245> A_IWL<6244> A_IWL<6243> A_IWL<6242> A_IWL<6241> A_IWL<6240> A_IWL<6239> A_IWL<6238> A_IWL<6237> A_IWL<6236> A_IWL<6235> A_IWL<6234> A_IWL<6233> A_IWL<6232> A_IWL<6231> A_IWL<6230> A_IWL<6229> A_IWL<6228> A_IWL<6227> A_IWL<6226> A_IWL<6225> A_IWL<6224> A_IWL<6223> A_IWL<6222> A_IWL<6221> A_IWL<6220> A_IWL<6219> A_IWL<6218> A_IWL<6217> A_IWL<6216> A_IWL<6215> A_IWL<6214> A_IWL<6213> A_IWL<6212> A_IWL<6211> A_IWL<6210> A_IWL<6209> A_IWL<6208> A_IWL<6207> A_IWL<6206> A_IWL<6205> A_IWL<6204> A_IWL<6203> A_IWL<6202> A_IWL<6201> A_IWL<6200> A_IWL<6199> A_IWL<6198> A_IWL<6197> A_IWL<6196> A_IWL<6195> A_IWL<6194> A_IWL<6193> A_IWL<6192> A_IWL<6191> A_IWL<6190> A_IWL<6189> A_IWL<6188> A_IWL<6187> A_IWL<6186> A_IWL<6185> A_IWL<6184> A_IWL<6183> A_IWL<6182> A_IWL<6181> A_IWL<6180> A_IWL<6179> A_IWL<6178> A_IWL<6177> A_IWL<6176> A_IWL<6175> A_IWL<6174> A_IWL<6173> A_IWL<6172> A_IWL<6171> A_IWL<6170> A_IWL<6169> A_IWL<6168> A_IWL<6167> A_IWL<6166> A_IWL<6165> A_IWL<6164> A_IWL<6163> A_IWL<6162> A_IWL<6161> A_IWL<6160> A_IWL<6159> A_IWL<6158> A_IWL<6157> A_IWL<6156> A_IWL<6155> A_IWL<6154> A_IWL<6153> A_IWL<6152> A_IWL<6151> A_IWL<6150> A_IWL<6149> A_IWL<6148> A_IWL<6147> A_IWL<6146> A_IWL<6145> A_IWL<6144> A_IWL<7167> A_IWL<7166> A_IWL<7165> A_IWL<7164> A_IWL<7163> A_IWL<7162> A_IWL<7161> A_IWL<7160> A_IWL<7159> A_IWL<7158> A_IWL<7157> A_IWL<7156> A_IWL<7155> A_IWL<7154> A_IWL<7153> A_IWL<7152> A_IWL<7151> A_IWL<7150> A_IWL<7149> A_IWL<7148> A_IWL<7147> A_IWL<7146> A_IWL<7145> A_IWL<7144> A_IWL<7143> A_IWL<7142> A_IWL<7141> A_IWL<7140> A_IWL<7139> A_IWL<7138> A_IWL<7137> A_IWL<7136> A_IWL<7135> A_IWL<7134> A_IWL<7133> A_IWL<7132> A_IWL<7131> A_IWL<7130> A_IWL<7129> A_IWL<7128> A_IWL<7127> A_IWL<7126> A_IWL<7125> A_IWL<7124> A_IWL<7123> A_IWL<7122> A_IWL<7121> A_IWL<7120> A_IWL<7119> A_IWL<7118> A_IWL<7117> A_IWL<7116> A_IWL<7115> A_IWL<7114> A_IWL<7113> A_IWL<7112> A_IWL<7111> A_IWL<7110> A_IWL<7109> A_IWL<7108> A_IWL<7107> A_IWL<7106> A_IWL<7105> A_IWL<7104> A_IWL<7103> A_IWL<7102> A_IWL<7101> A_IWL<7100> A_IWL<7099> A_IWL<7098> A_IWL<7097> A_IWL<7096> A_IWL<7095> A_IWL<7094> A_IWL<7093> A_IWL<7092> A_IWL<7091> A_IWL<7090> A_IWL<7089> A_IWL<7088> A_IWL<7087> A_IWL<7086> A_IWL<7085> A_IWL<7084> A_IWL<7083> A_IWL<7082> A_IWL<7081> A_IWL<7080> A_IWL<7079> A_IWL<7078> A_IWL<7077> A_IWL<7076> A_IWL<7075> A_IWL<7074> A_IWL<7073> A_IWL<7072> A_IWL<7071> A_IWL<7070> A_IWL<7069> A_IWL<7068> A_IWL<7067> A_IWL<7066> A_IWL<7065> A_IWL<7064> A_IWL<7063> A_IWL<7062> A_IWL<7061> A_IWL<7060> A_IWL<7059> A_IWL<7058> A_IWL<7057> A_IWL<7056> A_IWL<7055> A_IWL<7054> A_IWL<7053> A_IWL<7052> A_IWL<7051> A_IWL<7050> A_IWL<7049> A_IWL<7048> A_IWL<7047> A_IWL<7046> A_IWL<7045> A_IWL<7044> A_IWL<7043> A_IWL<7042> A_IWL<7041> A_IWL<7040> A_IWL<7039> A_IWL<7038> A_IWL<7037> A_IWL<7036> A_IWL<7035> A_IWL<7034> A_IWL<7033> A_IWL<7032> A_IWL<7031> A_IWL<7030> A_IWL<7029> A_IWL<7028> A_IWL<7027> A_IWL<7026> A_IWL<7025> A_IWL<7024> A_IWL<7023> A_IWL<7022> A_IWL<7021> A_IWL<7020> A_IWL<7019> A_IWL<7018> A_IWL<7017> A_IWL<7016> A_IWL<7015> A_IWL<7014> A_IWL<7013> A_IWL<7012> A_IWL<7011> A_IWL<7010> A_IWL<7009> A_IWL<7008> A_IWL<7007> A_IWL<7006> A_IWL<7005> A_IWL<7004> A_IWL<7003> A_IWL<7002> A_IWL<7001> A_IWL<7000> A_IWL<6999> A_IWL<6998> A_IWL<6997> A_IWL<6996> A_IWL<6995> A_IWL<6994> A_IWL<6993> A_IWL<6992> A_IWL<6991> A_IWL<6990> A_IWL<6989> A_IWL<6988> A_IWL<6987> A_IWL<6986> A_IWL<6985> A_IWL<6984> A_IWL<6983> A_IWL<6982> A_IWL<6981> A_IWL<6980> A_IWL<6979> A_IWL<6978> A_IWL<6977> A_IWL<6976> A_IWL<6975> A_IWL<6974> A_IWL<6973> A_IWL<6972> A_IWL<6971> A_IWL<6970> A_IWL<6969> A_IWL<6968> A_IWL<6967> A_IWL<6966> A_IWL<6965> A_IWL<6964> A_IWL<6963> A_IWL<6962> A_IWL<6961> A_IWL<6960> A_IWL<6959> A_IWL<6958> A_IWL<6957> A_IWL<6956> A_IWL<6955> A_IWL<6954> A_IWL<6953> A_IWL<6952> A_IWL<6951> A_IWL<6950> A_IWL<6949> A_IWL<6948> A_IWL<6947> A_IWL<6946> A_IWL<6945> A_IWL<6944> A_IWL<6943> A_IWL<6942> A_IWL<6941> A_IWL<6940> A_IWL<6939> A_IWL<6938> A_IWL<6937> A_IWL<6936> A_IWL<6935> A_IWL<6934> A_IWL<6933> A_IWL<6932> A_IWL<6931> A_IWL<6930> A_IWL<6929> A_IWL<6928> A_IWL<6927> A_IWL<6926> A_IWL<6925> A_IWL<6924> A_IWL<6923> A_IWL<6922> A_IWL<6921> A_IWL<6920> A_IWL<6919> A_IWL<6918> A_IWL<6917> A_IWL<6916> A_IWL<6915> A_IWL<6914> A_IWL<6913> A_IWL<6912> A_IWL<6911> A_IWL<6910> A_IWL<6909> A_IWL<6908> A_IWL<6907> A_IWL<6906> A_IWL<6905> A_IWL<6904> A_IWL<6903> A_IWL<6902> A_IWL<6901> A_IWL<6900> A_IWL<6899> A_IWL<6898> A_IWL<6897> A_IWL<6896> A_IWL<6895> A_IWL<6894> A_IWL<6893> A_IWL<6892> A_IWL<6891> A_IWL<6890> A_IWL<6889> A_IWL<6888> A_IWL<6887> A_IWL<6886> A_IWL<6885> A_IWL<6884> A_IWL<6883> A_IWL<6882> A_IWL<6881> A_IWL<6880> A_IWL<6879> A_IWL<6878> A_IWL<6877> A_IWL<6876> A_IWL<6875> A_IWL<6874> A_IWL<6873> A_IWL<6872> A_IWL<6871> A_IWL<6870> A_IWL<6869> A_IWL<6868> A_IWL<6867> A_IWL<6866> A_IWL<6865> A_IWL<6864> A_IWL<6863> A_IWL<6862> A_IWL<6861> A_IWL<6860> A_IWL<6859> A_IWL<6858> A_IWL<6857> A_IWL<6856> A_IWL<6855> A_IWL<6854> A_IWL<6853> A_IWL<6852> A_IWL<6851> A_IWL<6850> A_IWL<6849> A_IWL<6848> A_IWL<6847> A_IWL<6846> A_IWL<6845> A_IWL<6844> A_IWL<6843> A_IWL<6842> A_IWL<6841> A_IWL<6840> A_IWL<6839> A_IWL<6838> A_IWL<6837> A_IWL<6836> A_IWL<6835> A_IWL<6834> A_IWL<6833> A_IWL<6832> A_IWL<6831> A_IWL<6830> A_IWL<6829> A_IWL<6828> A_IWL<6827> A_IWL<6826> A_IWL<6825> A_IWL<6824> A_IWL<6823> A_IWL<6822> A_IWL<6821> A_IWL<6820> A_IWL<6819> A_IWL<6818> A_IWL<6817> A_IWL<6816> A_IWL<6815> A_IWL<6814> A_IWL<6813> A_IWL<6812> A_IWL<6811> A_IWL<6810> A_IWL<6809> A_IWL<6808> A_IWL<6807> A_IWL<6806> A_IWL<6805> A_IWL<6804> A_IWL<6803> A_IWL<6802> A_IWL<6801> A_IWL<6800> A_IWL<6799> A_IWL<6798> A_IWL<6797> A_IWL<6796> A_IWL<6795> A_IWL<6794> A_IWL<6793> A_IWL<6792> A_IWL<6791> A_IWL<6790> A_IWL<6789> A_IWL<6788> A_IWL<6787> A_IWL<6786> A_IWL<6785> A_IWL<6784> A_IWL<6783> A_IWL<6782> A_IWL<6781> A_IWL<6780> A_IWL<6779> A_IWL<6778> A_IWL<6777> A_IWL<6776> A_IWL<6775> A_IWL<6774> A_IWL<6773> A_IWL<6772> A_IWL<6771> A_IWL<6770> A_IWL<6769> A_IWL<6768> A_IWL<6767> A_IWL<6766> A_IWL<6765> A_IWL<6764> A_IWL<6763> A_IWL<6762> A_IWL<6761> A_IWL<6760> A_IWL<6759> A_IWL<6758> A_IWL<6757> A_IWL<6756> A_IWL<6755> A_IWL<6754> A_IWL<6753> A_IWL<6752> A_IWL<6751> A_IWL<6750> A_IWL<6749> A_IWL<6748> A_IWL<6747> A_IWL<6746> A_IWL<6745> A_IWL<6744> A_IWL<6743> A_IWL<6742> A_IWL<6741> A_IWL<6740> A_IWL<6739> A_IWL<6738> A_IWL<6737> A_IWL<6736> A_IWL<6735> A_IWL<6734> A_IWL<6733> A_IWL<6732> A_IWL<6731> A_IWL<6730> A_IWL<6729> A_IWL<6728> A_IWL<6727> A_IWL<6726> A_IWL<6725> A_IWL<6724> A_IWL<6723> A_IWL<6722> A_IWL<6721> A_IWL<6720> A_IWL<6719> A_IWL<6718> A_IWL<6717> A_IWL<6716> A_IWL<6715> A_IWL<6714> A_IWL<6713> A_IWL<6712> A_IWL<6711> A_IWL<6710> A_IWL<6709> A_IWL<6708> A_IWL<6707> A_IWL<6706> A_IWL<6705> A_IWL<6704> A_IWL<6703> A_IWL<6702> A_IWL<6701> A_IWL<6700> A_IWL<6699> A_IWL<6698> A_IWL<6697> A_IWL<6696> A_IWL<6695> A_IWL<6694> A_IWL<6693> A_IWL<6692> A_IWL<6691> A_IWL<6690> A_IWL<6689> A_IWL<6688> A_IWL<6687> A_IWL<6686> A_IWL<6685> A_IWL<6684> A_IWL<6683> A_IWL<6682> A_IWL<6681> A_IWL<6680> A_IWL<6679> A_IWL<6678> A_IWL<6677> A_IWL<6676> A_IWL<6675> A_IWL<6674> A_IWL<6673> A_IWL<6672> A_IWL<6671> A_IWL<6670> A_IWL<6669> A_IWL<6668> A_IWL<6667> A_IWL<6666> A_IWL<6665> A_IWL<6664> A_IWL<6663> A_IWL<6662> A_IWL<6661> A_IWL<6660> A_IWL<6659> A_IWL<6658> A_IWL<6657> A_IWL<6656> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<12> A_BLC<25> A_BLC<24> A_BLC_TOP<25> A_BLC_TOP<24> A_BLT<25> A_BLT<24> A_BLT_TOP<25> A_BLT_TOP<24> A_IWL<6143> A_IWL<6142> A_IWL<6141> A_IWL<6140> A_IWL<6139> A_IWL<6138> A_IWL<6137> A_IWL<6136> A_IWL<6135> A_IWL<6134> A_IWL<6133> A_IWL<6132> A_IWL<6131> A_IWL<6130> A_IWL<6129> A_IWL<6128> A_IWL<6127> A_IWL<6126> A_IWL<6125> A_IWL<6124> A_IWL<6123> A_IWL<6122> A_IWL<6121> A_IWL<6120> A_IWL<6119> A_IWL<6118> A_IWL<6117> A_IWL<6116> A_IWL<6115> A_IWL<6114> A_IWL<6113> A_IWL<6112> A_IWL<6111> A_IWL<6110> A_IWL<6109> A_IWL<6108> A_IWL<6107> A_IWL<6106> A_IWL<6105> A_IWL<6104> A_IWL<6103> A_IWL<6102> A_IWL<6101> A_IWL<6100> A_IWL<6099> A_IWL<6098> A_IWL<6097> A_IWL<6096> A_IWL<6095> A_IWL<6094> A_IWL<6093> A_IWL<6092> A_IWL<6091> A_IWL<6090> A_IWL<6089> A_IWL<6088> A_IWL<6087> A_IWL<6086> A_IWL<6085> A_IWL<6084> A_IWL<6083> A_IWL<6082> A_IWL<6081> A_IWL<6080> A_IWL<6079> A_IWL<6078> A_IWL<6077> A_IWL<6076> A_IWL<6075> A_IWL<6074> A_IWL<6073> A_IWL<6072> A_IWL<6071> A_IWL<6070> A_IWL<6069> A_IWL<6068> A_IWL<6067> A_IWL<6066> A_IWL<6065> A_IWL<6064> A_IWL<6063> A_IWL<6062> A_IWL<6061> A_IWL<6060> A_IWL<6059> A_IWL<6058> A_IWL<6057> A_IWL<6056> A_IWL<6055> A_IWL<6054> A_IWL<6053> A_IWL<6052> A_IWL<6051> A_IWL<6050> A_IWL<6049> A_IWL<6048> A_IWL<6047> A_IWL<6046> A_IWL<6045> A_IWL<6044> A_IWL<6043> A_IWL<6042> A_IWL<6041> A_IWL<6040> A_IWL<6039> A_IWL<6038> A_IWL<6037> A_IWL<6036> A_IWL<6035> A_IWL<6034> A_IWL<6033> A_IWL<6032> A_IWL<6031> A_IWL<6030> A_IWL<6029> A_IWL<6028> A_IWL<6027> A_IWL<6026> A_IWL<6025> A_IWL<6024> A_IWL<6023> A_IWL<6022> A_IWL<6021> A_IWL<6020> A_IWL<6019> A_IWL<6018> A_IWL<6017> A_IWL<6016> A_IWL<6015> A_IWL<6014> A_IWL<6013> A_IWL<6012> A_IWL<6011> A_IWL<6010> A_IWL<6009> A_IWL<6008> A_IWL<6007> A_IWL<6006> A_IWL<6005> A_IWL<6004> A_IWL<6003> A_IWL<6002> A_IWL<6001> A_IWL<6000> A_IWL<5999> A_IWL<5998> A_IWL<5997> A_IWL<5996> A_IWL<5995> A_IWL<5994> A_IWL<5993> A_IWL<5992> A_IWL<5991> A_IWL<5990> A_IWL<5989> A_IWL<5988> A_IWL<5987> A_IWL<5986> A_IWL<5985> A_IWL<5984> A_IWL<5983> A_IWL<5982> A_IWL<5981> A_IWL<5980> A_IWL<5979> A_IWL<5978> A_IWL<5977> A_IWL<5976> A_IWL<5975> A_IWL<5974> A_IWL<5973> A_IWL<5972> A_IWL<5971> A_IWL<5970> A_IWL<5969> A_IWL<5968> A_IWL<5967> A_IWL<5966> A_IWL<5965> A_IWL<5964> A_IWL<5963> A_IWL<5962> A_IWL<5961> A_IWL<5960> A_IWL<5959> A_IWL<5958> A_IWL<5957> A_IWL<5956> A_IWL<5955> A_IWL<5954> A_IWL<5953> A_IWL<5952> A_IWL<5951> A_IWL<5950> A_IWL<5949> A_IWL<5948> A_IWL<5947> A_IWL<5946> A_IWL<5945> A_IWL<5944> A_IWL<5943> A_IWL<5942> A_IWL<5941> A_IWL<5940> A_IWL<5939> A_IWL<5938> A_IWL<5937> A_IWL<5936> A_IWL<5935> A_IWL<5934> A_IWL<5933> A_IWL<5932> A_IWL<5931> A_IWL<5930> A_IWL<5929> A_IWL<5928> A_IWL<5927> A_IWL<5926> A_IWL<5925> A_IWL<5924> A_IWL<5923> A_IWL<5922> A_IWL<5921> A_IWL<5920> A_IWL<5919> A_IWL<5918> A_IWL<5917> A_IWL<5916> A_IWL<5915> A_IWL<5914> A_IWL<5913> A_IWL<5912> A_IWL<5911> A_IWL<5910> A_IWL<5909> A_IWL<5908> A_IWL<5907> A_IWL<5906> A_IWL<5905> A_IWL<5904> A_IWL<5903> A_IWL<5902> A_IWL<5901> A_IWL<5900> A_IWL<5899> A_IWL<5898> A_IWL<5897> A_IWL<5896> A_IWL<5895> A_IWL<5894> A_IWL<5893> A_IWL<5892> A_IWL<5891> A_IWL<5890> A_IWL<5889> A_IWL<5888> A_IWL<5887> A_IWL<5886> A_IWL<5885> A_IWL<5884> A_IWL<5883> A_IWL<5882> A_IWL<5881> A_IWL<5880> A_IWL<5879> A_IWL<5878> A_IWL<5877> A_IWL<5876> A_IWL<5875> A_IWL<5874> A_IWL<5873> A_IWL<5872> A_IWL<5871> A_IWL<5870> A_IWL<5869> A_IWL<5868> A_IWL<5867> A_IWL<5866> A_IWL<5865> A_IWL<5864> A_IWL<5863> A_IWL<5862> A_IWL<5861> A_IWL<5860> A_IWL<5859> A_IWL<5858> A_IWL<5857> A_IWL<5856> A_IWL<5855> A_IWL<5854> A_IWL<5853> A_IWL<5852> A_IWL<5851> A_IWL<5850> A_IWL<5849> A_IWL<5848> A_IWL<5847> A_IWL<5846> A_IWL<5845> A_IWL<5844> A_IWL<5843> A_IWL<5842> A_IWL<5841> A_IWL<5840> A_IWL<5839> A_IWL<5838> A_IWL<5837> A_IWL<5836> A_IWL<5835> A_IWL<5834> A_IWL<5833> A_IWL<5832> A_IWL<5831> A_IWL<5830> A_IWL<5829> A_IWL<5828> A_IWL<5827> A_IWL<5826> A_IWL<5825> A_IWL<5824> A_IWL<5823> A_IWL<5822> A_IWL<5821> A_IWL<5820> A_IWL<5819> A_IWL<5818> A_IWL<5817> A_IWL<5816> A_IWL<5815> A_IWL<5814> A_IWL<5813> A_IWL<5812> A_IWL<5811> A_IWL<5810> A_IWL<5809> A_IWL<5808> A_IWL<5807> A_IWL<5806> A_IWL<5805> A_IWL<5804> A_IWL<5803> A_IWL<5802> A_IWL<5801> A_IWL<5800> A_IWL<5799> A_IWL<5798> A_IWL<5797> A_IWL<5796> A_IWL<5795> A_IWL<5794> A_IWL<5793> A_IWL<5792> A_IWL<5791> A_IWL<5790> A_IWL<5789> A_IWL<5788> A_IWL<5787> A_IWL<5786> A_IWL<5785> A_IWL<5784> A_IWL<5783> A_IWL<5782> A_IWL<5781> A_IWL<5780> A_IWL<5779> A_IWL<5778> A_IWL<5777> A_IWL<5776> A_IWL<5775> A_IWL<5774> A_IWL<5773> A_IWL<5772> A_IWL<5771> A_IWL<5770> A_IWL<5769> A_IWL<5768> A_IWL<5767> A_IWL<5766> A_IWL<5765> A_IWL<5764> A_IWL<5763> A_IWL<5762> A_IWL<5761> A_IWL<5760> A_IWL<5759> A_IWL<5758> A_IWL<5757> A_IWL<5756> A_IWL<5755> A_IWL<5754> A_IWL<5753> A_IWL<5752> A_IWL<5751> A_IWL<5750> A_IWL<5749> A_IWL<5748> A_IWL<5747> A_IWL<5746> A_IWL<5745> A_IWL<5744> A_IWL<5743> A_IWL<5742> A_IWL<5741> A_IWL<5740> A_IWL<5739> A_IWL<5738> A_IWL<5737> A_IWL<5736> A_IWL<5735> A_IWL<5734> A_IWL<5733> A_IWL<5732> A_IWL<5731> A_IWL<5730> A_IWL<5729> A_IWL<5728> A_IWL<5727> A_IWL<5726> A_IWL<5725> A_IWL<5724> A_IWL<5723> A_IWL<5722> A_IWL<5721> A_IWL<5720> A_IWL<5719> A_IWL<5718> A_IWL<5717> A_IWL<5716> A_IWL<5715> A_IWL<5714> A_IWL<5713> A_IWL<5712> A_IWL<5711> A_IWL<5710> A_IWL<5709> A_IWL<5708> A_IWL<5707> A_IWL<5706> A_IWL<5705> A_IWL<5704> A_IWL<5703> A_IWL<5702> A_IWL<5701> A_IWL<5700> A_IWL<5699> A_IWL<5698> A_IWL<5697> A_IWL<5696> A_IWL<5695> A_IWL<5694> A_IWL<5693> A_IWL<5692> A_IWL<5691> A_IWL<5690> A_IWL<5689> A_IWL<5688> A_IWL<5687> A_IWL<5686> A_IWL<5685> A_IWL<5684> A_IWL<5683> A_IWL<5682> A_IWL<5681> A_IWL<5680> A_IWL<5679> A_IWL<5678> A_IWL<5677> A_IWL<5676> A_IWL<5675> A_IWL<5674> A_IWL<5673> A_IWL<5672> A_IWL<5671> A_IWL<5670> A_IWL<5669> A_IWL<5668> A_IWL<5667> A_IWL<5666> A_IWL<5665> A_IWL<5664> A_IWL<5663> A_IWL<5662> A_IWL<5661> A_IWL<5660> A_IWL<5659> A_IWL<5658> A_IWL<5657> A_IWL<5656> A_IWL<5655> A_IWL<5654> A_IWL<5653> A_IWL<5652> A_IWL<5651> A_IWL<5650> A_IWL<5649> A_IWL<5648> A_IWL<5647> A_IWL<5646> A_IWL<5645> A_IWL<5644> A_IWL<5643> A_IWL<5642> A_IWL<5641> A_IWL<5640> A_IWL<5639> A_IWL<5638> A_IWL<5637> A_IWL<5636> A_IWL<5635> A_IWL<5634> A_IWL<5633> A_IWL<5632> A_IWL<6655> A_IWL<6654> A_IWL<6653> A_IWL<6652> A_IWL<6651> A_IWL<6650> A_IWL<6649> A_IWL<6648> A_IWL<6647> A_IWL<6646> A_IWL<6645> A_IWL<6644> A_IWL<6643> A_IWL<6642> A_IWL<6641> A_IWL<6640> A_IWL<6639> A_IWL<6638> A_IWL<6637> A_IWL<6636> A_IWL<6635> A_IWL<6634> A_IWL<6633> A_IWL<6632> A_IWL<6631> A_IWL<6630> A_IWL<6629> A_IWL<6628> A_IWL<6627> A_IWL<6626> A_IWL<6625> A_IWL<6624> A_IWL<6623> A_IWL<6622> A_IWL<6621> A_IWL<6620> A_IWL<6619> A_IWL<6618> A_IWL<6617> A_IWL<6616> A_IWL<6615> A_IWL<6614> A_IWL<6613> A_IWL<6612> A_IWL<6611> A_IWL<6610> A_IWL<6609> A_IWL<6608> A_IWL<6607> A_IWL<6606> A_IWL<6605> A_IWL<6604> A_IWL<6603> A_IWL<6602> A_IWL<6601> A_IWL<6600> A_IWL<6599> A_IWL<6598> A_IWL<6597> A_IWL<6596> A_IWL<6595> A_IWL<6594> A_IWL<6593> A_IWL<6592> A_IWL<6591> A_IWL<6590> A_IWL<6589> A_IWL<6588> A_IWL<6587> A_IWL<6586> A_IWL<6585> A_IWL<6584> A_IWL<6583> A_IWL<6582> A_IWL<6581> A_IWL<6580> A_IWL<6579> A_IWL<6578> A_IWL<6577> A_IWL<6576> A_IWL<6575> A_IWL<6574> A_IWL<6573> A_IWL<6572> A_IWL<6571> A_IWL<6570> A_IWL<6569> A_IWL<6568> A_IWL<6567> A_IWL<6566> A_IWL<6565> A_IWL<6564> A_IWL<6563> A_IWL<6562> A_IWL<6561> A_IWL<6560> A_IWL<6559> A_IWL<6558> A_IWL<6557> A_IWL<6556> A_IWL<6555> A_IWL<6554> A_IWL<6553> A_IWL<6552> A_IWL<6551> A_IWL<6550> A_IWL<6549> A_IWL<6548> A_IWL<6547> A_IWL<6546> A_IWL<6545> A_IWL<6544> A_IWL<6543> A_IWL<6542> A_IWL<6541> A_IWL<6540> A_IWL<6539> A_IWL<6538> A_IWL<6537> A_IWL<6536> A_IWL<6535> A_IWL<6534> A_IWL<6533> A_IWL<6532> A_IWL<6531> A_IWL<6530> A_IWL<6529> A_IWL<6528> A_IWL<6527> A_IWL<6526> A_IWL<6525> A_IWL<6524> A_IWL<6523> A_IWL<6522> A_IWL<6521> A_IWL<6520> A_IWL<6519> A_IWL<6518> A_IWL<6517> A_IWL<6516> A_IWL<6515> A_IWL<6514> A_IWL<6513> A_IWL<6512> A_IWL<6511> A_IWL<6510> A_IWL<6509> A_IWL<6508> A_IWL<6507> A_IWL<6506> A_IWL<6505> A_IWL<6504> A_IWL<6503> A_IWL<6502> A_IWL<6501> A_IWL<6500> A_IWL<6499> A_IWL<6498> A_IWL<6497> A_IWL<6496> A_IWL<6495> A_IWL<6494> A_IWL<6493> A_IWL<6492> A_IWL<6491> A_IWL<6490> A_IWL<6489> A_IWL<6488> A_IWL<6487> A_IWL<6486> A_IWL<6485> A_IWL<6484> A_IWL<6483> A_IWL<6482> A_IWL<6481> A_IWL<6480> A_IWL<6479> A_IWL<6478> A_IWL<6477> A_IWL<6476> A_IWL<6475> A_IWL<6474> A_IWL<6473> A_IWL<6472> A_IWL<6471> A_IWL<6470> A_IWL<6469> A_IWL<6468> A_IWL<6467> A_IWL<6466> A_IWL<6465> A_IWL<6464> A_IWL<6463> A_IWL<6462> A_IWL<6461> A_IWL<6460> A_IWL<6459> A_IWL<6458> A_IWL<6457> A_IWL<6456> A_IWL<6455> A_IWL<6454> A_IWL<6453> A_IWL<6452> A_IWL<6451> A_IWL<6450> A_IWL<6449> A_IWL<6448> A_IWL<6447> A_IWL<6446> A_IWL<6445> A_IWL<6444> A_IWL<6443> A_IWL<6442> A_IWL<6441> A_IWL<6440> A_IWL<6439> A_IWL<6438> A_IWL<6437> A_IWL<6436> A_IWL<6435> A_IWL<6434> A_IWL<6433> A_IWL<6432> A_IWL<6431> A_IWL<6430> A_IWL<6429> A_IWL<6428> A_IWL<6427> A_IWL<6426> A_IWL<6425> A_IWL<6424> A_IWL<6423> A_IWL<6422> A_IWL<6421> A_IWL<6420> A_IWL<6419> A_IWL<6418> A_IWL<6417> A_IWL<6416> A_IWL<6415> A_IWL<6414> A_IWL<6413> A_IWL<6412> A_IWL<6411> A_IWL<6410> A_IWL<6409> A_IWL<6408> A_IWL<6407> A_IWL<6406> A_IWL<6405> A_IWL<6404> A_IWL<6403> A_IWL<6402> A_IWL<6401> A_IWL<6400> A_IWL<6399> A_IWL<6398> A_IWL<6397> A_IWL<6396> A_IWL<6395> A_IWL<6394> A_IWL<6393> A_IWL<6392> A_IWL<6391> A_IWL<6390> A_IWL<6389> A_IWL<6388> A_IWL<6387> A_IWL<6386> A_IWL<6385> A_IWL<6384> A_IWL<6383> A_IWL<6382> A_IWL<6381> A_IWL<6380> A_IWL<6379> A_IWL<6378> A_IWL<6377> A_IWL<6376> A_IWL<6375> A_IWL<6374> A_IWL<6373> A_IWL<6372> A_IWL<6371> A_IWL<6370> A_IWL<6369> A_IWL<6368> A_IWL<6367> A_IWL<6366> A_IWL<6365> A_IWL<6364> A_IWL<6363> A_IWL<6362> A_IWL<6361> A_IWL<6360> A_IWL<6359> A_IWL<6358> A_IWL<6357> A_IWL<6356> A_IWL<6355> A_IWL<6354> A_IWL<6353> A_IWL<6352> A_IWL<6351> A_IWL<6350> A_IWL<6349> A_IWL<6348> A_IWL<6347> A_IWL<6346> A_IWL<6345> A_IWL<6344> A_IWL<6343> A_IWL<6342> A_IWL<6341> A_IWL<6340> A_IWL<6339> A_IWL<6338> A_IWL<6337> A_IWL<6336> A_IWL<6335> A_IWL<6334> A_IWL<6333> A_IWL<6332> A_IWL<6331> A_IWL<6330> A_IWL<6329> A_IWL<6328> A_IWL<6327> A_IWL<6326> A_IWL<6325> A_IWL<6324> A_IWL<6323> A_IWL<6322> A_IWL<6321> A_IWL<6320> A_IWL<6319> A_IWL<6318> A_IWL<6317> A_IWL<6316> A_IWL<6315> A_IWL<6314> A_IWL<6313> A_IWL<6312> A_IWL<6311> A_IWL<6310> A_IWL<6309> A_IWL<6308> A_IWL<6307> A_IWL<6306> A_IWL<6305> A_IWL<6304> A_IWL<6303> A_IWL<6302> A_IWL<6301> A_IWL<6300> A_IWL<6299> A_IWL<6298> A_IWL<6297> A_IWL<6296> A_IWL<6295> A_IWL<6294> A_IWL<6293> A_IWL<6292> A_IWL<6291> A_IWL<6290> A_IWL<6289> A_IWL<6288> A_IWL<6287> A_IWL<6286> A_IWL<6285> A_IWL<6284> A_IWL<6283> A_IWL<6282> A_IWL<6281> A_IWL<6280> A_IWL<6279> A_IWL<6278> A_IWL<6277> A_IWL<6276> A_IWL<6275> A_IWL<6274> A_IWL<6273> A_IWL<6272> A_IWL<6271> A_IWL<6270> A_IWL<6269> A_IWL<6268> A_IWL<6267> A_IWL<6266> A_IWL<6265> A_IWL<6264> A_IWL<6263> A_IWL<6262> A_IWL<6261> A_IWL<6260> A_IWL<6259> A_IWL<6258> A_IWL<6257> A_IWL<6256> A_IWL<6255> A_IWL<6254> A_IWL<6253> A_IWL<6252> A_IWL<6251> A_IWL<6250> A_IWL<6249> A_IWL<6248> A_IWL<6247> A_IWL<6246> A_IWL<6245> A_IWL<6244> A_IWL<6243> A_IWL<6242> A_IWL<6241> A_IWL<6240> A_IWL<6239> A_IWL<6238> A_IWL<6237> A_IWL<6236> A_IWL<6235> A_IWL<6234> A_IWL<6233> A_IWL<6232> A_IWL<6231> A_IWL<6230> A_IWL<6229> A_IWL<6228> A_IWL<6227> A_IWL<6226> A_IWL<6225> A_IWL<6224> A_IWL<6223> A_IWL<6222> A_IWL<6221> A_IWL<6220> A_IWL<6219> A_IWL<6218> A_IWL<6217> A_IWL<6216> A_IWL<6215> A_IWL<6214> A_IWL<6213> A_IWL<6212> A_IWL<6211> A_IWL<6210> A_IWL<6209> A_IWL<6208> A_IWL<6207> A_IWL<6206> A_IWL<6205> A_IWL<6204> A_IWL<6203> A_IWL<6202> A_IWL<6201> A_IWL<6200> A_IWL<6199> A_IWL<6198> A_IWL<6197> A_IWL<6196> A_IWL<6195> A_IWL<6194> A_IWL<6193> A_IWL<6192> A_IWL<6191> A_IWL<6190> A_IWL<6189> A_IWL<6188> A_IWL<6187> A_IWL<6186> A_IWL<6185> A_IWL<6184> A_IWL<6183> A_IWL<6182> A_IWL<6181> A_IWL<6180> A_IWL<6179> A_IWL<6178> A_IWL<6177> A_IWL<6176> A_IWL<6175> A_IWL<6174> A_IWL<6173> A_IWL<6172> A_IWL<6171> A_IWL<6170> A_IWL<6169> A_IWL<6168> A_IWL<6167> A_IWL<6166> A_IWL<6165> A_IWL<6164> A_IWL<6163> A_IWL<6162> A_IWL<6161> A_IWL<6160> A_IWL<6159> A_IWL<6158> A_IWL<6157> A_IWL<6156> A_IWL<6155> A_IWL<6154> A_IWL<6153> A_IWL<6152> A_IWL<6151> A_IWL<6150> A_IWL<6149> A_IWL<6148> A_IWL<6147> A_IWL<6146> A_IWL<6145> A_IWL<6144> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<11> A_BLC<23> A_BLC<22> A_BLC_TOP<23> A_BLC_TOP<22> A_BLT<23> A_BLT<22> A_BLT_TOP<23> A_BLT_TOP<22> A_IWL<5631> A_IWL<5630> A_IWL<5629> A_IWL<5628> A_IWL<5627> A_IWL<5626> A_IWL<5625> A_IWL<5624> A_IWL<5623> A_IWL<5622> A_IWL<5621> A_IWL<5620> A_IWL<5619> A_IWL<5618> A_IWL<5617> A_IWL<5616> A_IWL<5615> A_IWL<5614> A_IWL<5613> A_IWL<5612> A_IWL<5611> A_IWL<5610> A_IWL<5609> A_IWL<5608> A_IWL<5607> A_IWL<5606> A_IWL<5605> A_IWL<5604> A_IWL<5603> A_IWL<5602> A_IWL<5601> A_IWL<5600> A_IWL<5599> A_IWL<5598> A_IWL<5597> A_IWL<5596> A_IWL<5595> A_IWL<5594> A_IWL<5593> A_IWL<5592> A_IWL<5591> A_IWL<5590> A_IWL<5589> A_IWL<5588> A_IWL<5587> A_IWL<5586> A_IWL<5585> A_IWL<5584> A_IWL<5583> A_IWL<5582> A_IWL<5581> A_IWL<5580> A_IWL<5579> A_IWL<5578> A_IWL<5577> A_IWL<5576> A_IWL<5575> A_IWL<5574> A_IWL<5573> A_IWL<5572> A_IWL<5571> A_IWL<5570> A_IWL<5569> A_IWL<5568> A_IWL<5567> A_IWL<5566> A_IWL<5565> A_IWL<5564> A_IWL<5563> A_IWL<5562> A_IWL<5561> A_IWL<5560> A_IWL<5559> A_IWL<5558> A_IWL<5557> A_IWL<5556> A_IWL<5555> A_IWL<5554> A_IWL<5553> A_IWL<5552> A_IWL<5551> A_IWL<5550> A_IWL<5549> A_IWL<5548> A_IWL<5547> A_IWL<5546> A_IWL<5545> A_IWL<5544> A_IWL<5543> A_IWL<5542> A_IWL<5541> A_IWL<5540> A_IWL<5539> A_IWL<5538> A_IWL<5537> A_IWL<5536> A_IWL<5535> A_IWL<5534> A_IWL<5533> A_IWL<5532> A_IWL<5531> A_IWL<5530> A_IWL<5529> A_IWL<5528> A_IWL<5527> A_IWL<5526> A_IWL<5525> A_IWL<5524> A_IWL<5523> A_IWL<5522> A_IWL<5521> A_IWL<5520> A_IWL<5519> A_IWL<5518> A_IWL<5517> A_IWL<5516> A_IWL<5515> A_IWL<5514> A_IWL<5513> A_IWL<5512> A_IWL<5511> A_IWL<5510> A_IWL<5509> A_IWL<5508> A_IWL<5507> A_IWL<5506> A_IWL<5505> A_IWL<5504> A_IWL<5503> A_IWL<5502> A_IWL<5501> A_IWL<5500> A_IWL<5499> A_IWL<5498> A_IWL<5497> A_IWL<5496> A_IWL<5495> A_IWL<5494> A_IWL<5493> A_IWL<5492> A_IWL<5491> A_IWL<5490> A_IWL<5489> A_IWL<5488> A_IWL<5487> A_IWL<5486> A_IWL<5485> A_IWL<5484> A_IWL<5483> A_IWL<5482> A_IWL<5481> A_IWL<5480> A_IWL<5479> A_IWL<5478> A_IWL<5477> A_IWL<5476> A_IWL<5475> A_IWL<5474> A_IWL<5473> A_IWL<5472> A_IWL<5471> A_IWL<5470> A_IWL<5469> A_IWL<5468> A_IWL<5467> A_IWL<5466> A_IWL<5465> A_IWL<5464> A_IWL<5463> A_IWL<5462> A_IWL<5461> A_IWL<5460> A_IWL<5459> A_IWL<5458> A_IWL<5457> A_IWL<5456> A_IWL<5455> A_IWL<5454> A_IWL<5453> A_IWL<5452> A_IWL<5451> A_IWL<5450> A_IWL<5449> A_IWL<5448> A_IWL<5447> A_IWL<5446> A_IWL<5445> A_IWL<5444> A_IWL<5443> A_IWL<5442> A_IWL<5441> A_IWL<5440> A_IWL<5439> A_IWL<5438> A_IWL<5437> A_IWL<5436> A_IWL<5435> A_IWL<5434> A_IWL<5433> A_IWL<5432> A_IWL<5431> A_IWL<5430> A_IWL<5429> A_IWL<5428> A_IWL<5427> A_IWL<5426> A_IWL<5425> A_IWL<5424> A_IWL<5423> A_IWL<5422> A_IWL<5421> A_IWL<5420> A_IWL<5419> A_IWL<5418> A_IWL<5417> A_IWL<5416> A_IWL<5415> A_IWL<5414> A_IWL<5413> A_IWL<5412> A_IWL<5411> A_IWL<5410> A_IWL<5409> A_IWL<5408> A_IWL<5407> A_IWL<5406> A_IWL<5405> A_IWL<5404> A_IWL<5403> A_IWL<5402> A_IWL<5401> A_IWL<5400> A_IWL<5399> A_IWL<5398> A_IWL<5397> A_IWL<5396> A_IWL<5395> A_IWL<5394> A_IWL<5393> A_IWL<5392> A_IWL<5391> A_IWL<5390> A_IWL<5389> A_IWL<5388> A_IWL<5387> A_IWL<5386> A_IWL<5385> A_IWL<5384> A_IWL<5383> A_IWL<5382> A_IWL<5381> A_IWL<5380> A_IWL<5379> A_IWL<5378> A_IWL<5377> A_IWL<5376> A_IWL<5375> A_IWL<5374> A_IWL<5373> A_IWL<5372> A_IWL<5371> A_IWL<5370> A_IWL<5369> A_IWL<5368> A_IWL<5367> A_IWL<5366> A_IWL<5365> A_IWL<5364> A_IWL<5363> A_IWL<5362> A_IWL<5361> A_IWL<5360> A_IWL<5359> A_IWL<5358> A_IWL<5357> A_IWL<5356> A_IWL<5355> A_IWL<5354> A_IWL<5353> A_IWL<5352> A_IWL<5351> A_IWL<5350> A_IWL<5349> A_IWL<5348> A_IWL<5347> A_IWL<5346> A_IWL<5345> A_IWL<5344> A_IWL<5343> A_IWL<5342> A_IWL<5341> A_IWL<5340> A_IWL<5339> A_IWL<5338> A_IWL<5337> A_IWL<5336> A_IWL<5335> A_IWL<5334> A_IWL<5333> A_IWL<5332> A_IWL<5331> A_IWL<5330> A_IWL<5329> A_IWL<5328> A_IWL<5327> A_IWL<5326> A_IWL<5325> A_IWL<5324> A_IWL<5323> A_IWL<5322> A_IWL<5321> A_IWL<5320> A_IWL<5319> A_IWL<5318> A_IWL<5317> A_IWL<5316> A_IWL<5315> A_IWL<5314> A_IWL<5313> A_IWL<5312> A_IWL<5311> A_IWL<5310> A_IWL<5309> A_IWL<5308> A_IWL<5307> A_IWL<5306> A_IWL<5305> A_IWL<5304> A_IWL<5303> A_IWL<5302> A_IWL<5301> A_IWL<5300> A_IWL<5299> A_IWL<5298> A_IWL<5297> A_IWL<5296> A_IWL<5295> A_IWL<5294> A_IWL<5293> A_IWL<5292> A_IWL<5291> A_IWL<5290> A_IWL<5289> A_IWL<5288> A_IWL<5287> A_IWL<5286> A_IWL<5285> A_IWL<5284> A_IWL<5283> A_IWL<5282> A_IWL<5281> A_IWL<5280> A_IWL<5279> A_IWL<5278> A_IWL<5277> A_IWL<5276> A_IWL<5275> A_IWL<5274> A_IWL<5273> A_IWL<5272> A_IWL<5271> A_IWL<5270> A_IWL<5269> A_IWL<5268> A_IWL<5267> A_IWL<5266> A_IWL<5265> A_IWL<5264> A_IWL<5263> A_IWL<5262> A_IWL<5261> A_IWL<5260> A_IWL<5259> A_IWL<5258> A_IWL<5257> A_IWL<5256> A_IWL<5255> A_IWL<5254> A_IWL<5253> A_IWL<5252> A_IWL<5251> A_IWL<5250> A_IWL<5249> A_IWL<5248> A_IWL<5247> A_IWL<5246> A_IWL<5245> A_IWL<5244> A_IWL<5243> A_IWL<5242> A_IWL<5241> A_IWL<5240> A_IWL<5239> A_IWL<5238> A_IWL<5237> A_IWL<5236> A_IWL<5235> A_IWL<5234> A_IWL<5233> A_IWL<5232> A_IWL<5231> A_IWL<5230> A_IWL<5229> A_IWL<5228> A_IWL<5227> A_IWL<5226> A_IWL<5225> A_IWL<5224> A_IWL<5223> A_IWL<5222> A_IWL<5221> A_IWL<5220> A_IWL<5219> A_IWL<5218> A_IWL<5217> A_IWL<5216> A_IWL<5215> A_IWL<5214> A_IWL<5213> A_IWL<5212> A_IWL<5211> A_IWL<5210> A_IWL<5209> A_IWL<5208> A_IWL<5207> A_IWL<5206> A_IWL<5205> A_IWL<5204> A_IWL<5203> A_IWL<5202> A_IWL<5201> A_IWL<5200> A_IWL<5199> A_IWL<5198> A_IWL<5197> A_IWL<5196> A_IWL<5195> A_IWL<5194> A_IWL<5193> A_IWL<5192> A_IWL<5191> A_IWL<5190> A_IWL<5189> A_IWL<5188> A_IWL<5187> A_IWL<5186> A_IWL<5185> A_IWL<5184> A_IWL<5183> A_IWL<5182> A_IWL<5181> A_IWL<5180> A_IWL<5179> A_IWL<5178> A_IWL<5177> A_IWL<5176> A_IWL<5175> A_IWL<5174> A_IWL<5173> A_IWL<5172> A_IWL<5171> A_IWL<5170> A_IWL<5169> A_IWL<5168> A_IWL<5167> A_IWL<5166> A_IWL<5165> A_IWL<5164> A_IWL<5163> A_IWL<5162> A_IWL<5161> A_IWL<5160> A_IWL<5159> A_IWL<5158> A_IWL<5157> A_IWL<5156> A_IWL<5155> A_IWL<5154> A_IWL<5153> A_IWL<5152> A_IWL<5151> A_IWL<5150> A_IWL<5149> A_IWL<5148> A_IWL<5147> A_IWL<5146> A_IWL<5145> A_IWL<5144> A_IWL<5143> A_IWL<5142> A_IWL<5141> A_IWL<5140> A_IWL<5139> A_IWL<5138> A_IWL<5137> A_IWL<5136> A_IWL<5135> A_IWL<5134> A_IWL<5133> A_IWL<5132> A_IWL<5131> A_IWL<5130> A_IWL<5129> A_IWL<5128> A_IWL<5127> A_IWL<5126> A_IWL<5125> A_IWL<5124> A_IWL<5123> A_IWL<5122> A_IWL<5121> A_IWL<5120> A_IWL<6143> A_IWL<6142> A_IWL<6141> A_IWL<6140> A_IWL<6139> A_IWL<6138> A_IWL<6137> A_IWL<6136> A_IWL<6135> A_IWL<6134> A_IWL<6133> A_IWL<6132> A_IWL<6131> A_IWL<6130> A_IWL<6129> A_IWL<6128> A_IWL<6127> A_IWL<6126> A_IWL<6125> A_IWL<6124> A_IWL<6123> A_IWL<6122> A_IWL<6121> A_IWL<6120> A_IWL<6119> A_IWL<6118> A_IWL<6117> A_IWL<6116> A_IWL<6115> A_IWL<6114> A_IWL<6113> A_IWL<6112> A_IWL<6111> A_IWL<6110> A_IWL<6109> A_IWL<6108> A_IWL<6107> A_IWL<6106> A_IWL<6105> A_IWL<6104> A_IWL<6103> A_IWL<6102> A_IWL<6101> A_IWL<6100> A_IWL<6099> A_IWL<6098> A_IWL<6097> A_IWL<6096> A_IWL<6095> A_IWL<6094> A_IWL<6093> A_IWL<6092> A_IWL<6091> A_IWL<6090> A_IWL<6089> A_IWL<6088> A_IWL<6087> A_IWL<6086> A_IWL<6085> A_IWL<6084> A_IWL<6083> A_IWL<6082> A_IWL<6081> A_IWL<6080> A_IWL<6079> A_IWL<6078> A_IWL<6077> A_IWL<6076> A_IWL<6075> A_IWL<6074> A_IWL<6073> A_IWL<6072> A_IWL<6071> A_IWL<6070> A_IWL<6069> A_IWL<6068> A_IWL<6067> A_IWL<6066> A_IWL<6065> A_IWL<6064> A_IWL<6063> A_IWL<6062> A_IWL<6061> A_IWL<6060> A_IWL<6059> A_IWL<6058> A_IWL<6057> A_IWL<6056> A_IWL<6055> A_IWL<6054> A_IWL<6053> A_IWL<6052> A_IWL<6051> A_IWL<6050> A_IWL<6049> A_IWL<6048> A_IWL<6047> A_IWL<6046> A_IWL<6045> A_IWL<6044> A_IWL<6043> A_IWL<6042> A_IWL<6041> A_IWL<6040> A_IWL<6039> A_IWL<6038> A_IWL<6037> A_IWL<6036> A_IWL<6035> A_IWL<6034> A_IWL<6033> A_IWL<6032> A_IWL<6031> A_IWL<6030> A_IWL<6029> A_IWL<6028> A_IWL<6027> A_IWL<6026> A_IWL<6025> A_IWL<6024> A_IWL<6023> A_IWL<6022> A_IWL<6021> A_IWL<6020> A_IWL<6019> A_IWL<6018> A_IWL<6017> A_IWL<6016> A_IWL<6015> A_IWL<6014> A_IWL<6013> A_IWL<6012> A_IWL<6011> A_IWL<6010> A_IWL<6009> A_IWL<6008> A_IWL<6007> A_IWL<6006> A_IWL<6005> A_IWL<6004> A_IWL<6003> A_IWL<6002> A_IWL<6001> A_IWL<6000> A_IWL<5999> A_IWL<5998> A_IWL<5997> A_IWL<5996> A_IWL<5995> A_IWL<5994> A_IWL<5993> A_IWL<5992> A_IWL<5991> A_IWL<5990> A_IWL<5989> A_IWL<5988> A_IWL<5987> A_IWL<5986> A_IWL<5985> A_IWL<5984> A_IWL<5983> A_IWL<5982> A_IWL<5981> A_IWL<5980> A_IWL<5979> A_IWL<5978> A_IWL<5977> A_IWL<5976> A_IWL<5975> A_IWL<5974> A_IWL<5973> A_IWL<5972> A_IWL<5971> A_IWL<5970> A_IWL<5969> A_IWL<5968> A_IWL<5967> A_IWL<5966> A_IWL<5965> A_IWL<5964> A_IWL<5963> A_IWL<5962> A_IWL<5961> A_IWL<5960> A_IWL<5959> A_IWL<5958> A_IWL<5957> A_IWL<5956> A_IWL<5955> A_IWL<5954> A_IWL<5953> A_IWL<5952> A_IWL<5951> A_IWL<5950> A_IWL<5949> A_IWL<5948> A_IWL<5947> A_IWL<5946> A_IWL<5945> A_IWL<5944> A_IWL<5943> A_IWL<5942> A_IWL<5941> A_IWL<5940> A_IWL<5939> A_IWL<5938> A_IWL<5937> A_IWL<5936> A_IWL<5935> A_IWL<5934> A_IWL<5933> A_IWL<5932> A_IWL<5931> A_IWL<5930> A_IWL<5929> A_IWL<5928> A_IWL<5927> A_IWL<5926> A_IWL<5925> A_IWL<5924> A_IWL<5923> A_IWL<5922> A_IWL<5921> A_IWL<5920> A_IWL<5919> A_IWL<5918> A_IWL<5917> A_IWL<5916> A_IWL<5915> A_IWL<5914> A_IWL<5913> A_IWL<5912> A_IWL<5911> A_IWL<5910> A_IWL<5909> A_IWL<5908> A_IWL<5907> A_IWL<5906> A_IWL<5905> A_IWL<5904> A_IWL<5903> A_IWL<5902> A_IWL<5901> A_IWL<5900> A_IWL<5899> A_IWL<5898> A_IWL<5897> A_IWL<5896> A_IWL<5895> A_IWL<5894> A_IWL<5893> A_IWL<5892> A_IWL<5891> A_IWL<5890> A_IWL<5889> A_IWL<5888> A_IWL<5887> A_IWL<5886> A_IWL<5885> A_IWL<5884> A_IWL<5883> A_IWL<5882> A_IWL<5881> A_IWL<5880> A_IWL<5879> A_IWL<5878> A_IWL<5877> A_IWL<5876> A_IWL<5875> A_IWL<5874> A_IWL<5873> A_IWL<5872> A_IWL<5871> A_IWL<5870> A_IWL<5869> A_IWL<5868> A_IWL<5867> A_IWL<5866> A_IWL<5865> A_IWL<5864> A_IWL<5863> A_IWL<5862> A_IWL<5861> A_IWL<5860> A_IWL<5859> A_IWL<5858> A_IWL<5857> A_IWL<5856> A_IWL<5855> A_IWL<5854> A_IWL<5853> A_IWL<5852> A_IWL<5851> A_IWL<5850> A_IWL<5849> A_IWL<5848> A_IWL<5847> A_IWL<5846> A_IWL<5845> A_IWL<5844> A_IWL<5843> A_IWL<5842> A_IWL<5841> A_IWL<5840> A_IWL<5839> A_IWL<5838> A_IWL<5837> A_IWL<5836> A_IWL<5835> A_IWL<5834> A_IWL<5833> A_IWL<5832> A_IWL<5831> A_IWL<5830> A_IWL<5829> A_IWL<5828> A_IWL<5827> A_IWL<5826> A_IWL<5825> A_IWL<5824> A_IWL<5823> A_IWL<5822> A_IWL<5821> A_IWL<5820> A_IWL<5819> A_IWL<5818> A_IWL<5817> A_IWL<5816> A_IWL<5815> A_IWL<5814> A_IWL<5813> A_IWL<5812> A_IWL<5811> A_IWL<5810> A_IWL<5809> A_IWL<5808> A_IWL<5807> A_IWL<5806> A_IWL<5805> A_IWL<5804> A_IWL<5803> A_IWL<5802> A_IWL<5801> A_IWL<5800> A_IWL<5799> A_IWL<5798> A_IWL<5797> A_IWL<5796> A_IWL<5795> A_IWL<5794> A_IWL<5793> A_IWL<5792> A_IWL<5791> A_IWL<5790> A_IWL<5789> A_IWL<5788> A_IWL<5787> A_IWL<5786> A_IWL<5785> A_IWL<5784> A_IWL<5783> A_IWL<5782> A_IWL<5781> A_IWL<5780> A_IWL<5779> A_IWL<5778> A_IWL<5777> A_IWL<5776> A_IWL<5775> A_IWL<5774> A_IWL<5773> A_IWL<5772> A_IWL<5771> A_IWL<5770> A_IWL<5769> A_IWL<5768> A_IWL<5767> A_IWL<5766> A_IWL<5765> A_IWL<5764> A_IWL<5763> A_IWL<5762> A_IWL<5761> A_IWL<5760> A_IWL<5759> A_IWL<5758> A_IWL<5757> A_IWL<5756> A_IWL<5755> A_IWL<5754> A_IWL<5753> A_IWL<5752> A_IWL<5751> A_IWL<5750> A_IWL<5749> A_IWL<5748> A_IWL<5747> A_IWL<5746> A_IWL<5745> A_IWL<5744> A_IWL<5743> A_IWL<5742> A_IWL<5741> A_IWL<5740> A_IWL<5739> A_IWL<5738> A_IWL<5737> A_IWL<5736> A_IWL<5735> A_IWL<5734> A_IWL<5733> A_IWL<5732> A_IWL<5731> A_IWL<5730> A_IWL<5729> A_IWL<5728> A_IWL<5727> A_IWL<5726> A_IWL<5725> A_IWL<5724> A_IWL<5723> A_IWL<5722> A_IWL<5721> A_IWL<5720> A_IWL<5719> A_IWL<5718> A_IWL<5717> A_IWL<5716> A_IWL<5715> A_IWL<5714> A_IWL<5713> A_IWL<5712> A_IWL<5711> A_IWL<5710> A_IWL<5709> A_IWL<5708> A_IWL<5707> A_IWL<5706> A_IWL<5705> A_IWL<5704> A_IWL<5703> A_IWL<5702> A_IWL<5701> A_IWL<5700> A_IWL<5699> A_IWL<5698> A_IWL<5697> A_IWL<5696> A_IWL<5695> A_IWL<5694> A_IWL<5693> A_IWL<5692> A_IWL<5691> A_IWL<5690> A_IWL<5689> A_IWL<5688> A_IWL<5687> A_IWL<5686> A_IWL<5685> A_IWL<5684> A_IWL<5683> A_IWL<5682> A_IWL<5681> A_IWL<5680> A_IWL<5679> A_IWL<5678> A_IWL<5677> A_IWL<5676> A_IWL<5675> A_IWL<5674> A_IWL<5673> A_IWL<5672> A_IWL<5671> A_IWL<5670> A_IWL<5669> A_IWL<5668> A_IWL<5667> A_IWL<5666> A_IWL<5665> A_IWL<5664> A_IWL<5663> A_IWL<5662> A_IWL<5661> A_IWL<5660> A_IWL<5659> A_IWL<5658> A_IWL<5657> A_IWL<5656> A_IWL<5655> A_IWL<5654> A_IWL<5653> A_IWL<5652> A_IWL<5651> A_IWL<5650> A_IWL<5649> A_IWL<5648> A_IWL<5647> A_IWL<5646> A_IWL<5645> A_IWL<5644> A_IWL<5643> A_IWL<5642> A_IWL<5641> A_IWL<5640> A_IWL<5639> A_IWL<5638> A_IWL<5637> A_IWL<5636> A_IWL<5635> A_IWL<5634> A_IWL<5633> A_IWL<5632> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<10> A_BLC<21> A_BLC<20> A_BLC_TOP<21> A_BLC_TOP<20> A_BLT<21> A_BLT<20> A_BLT_TOP<21> A_BLT_TOP<20> A_IWL<5119> A_IWL<5118> A_IWL<5117> A_IWL<5116> A_IWL<5115> A_IWL<5114> A_IWL<5113> A_IWL<5112> A_IWL<5111> A_IWL<5110> A_IWL<5109> A_IWL<5108> A_IWL<5107> A_IWL<5106> A_IWL<5105> A_IWL<5104> A_IWL<5103> A_IWL<5102> A_IWL<5101> A_IWL<5100> A_IWL<5099> A_IWL<5098> A_IWL<5097> A_IWL<5096> A_IWL<5095> A_IWL<5094> A_IWL<5093> A_IWL<5092> A_IWL<5091> A_IWL<5090> A_IWL<5089> A_IWL<5088> A_IWL<5087> A_IWL<5086> A_IWL<5085> A_IWL<5084> A_IWL<5083> A_IWL<5082> A_IWL<5081> A_IWL<5080> A_IWL<5079> A_IWL<5078> A_IWL<5077> A_IWL<5076> A_IWL<5075> A_IWL<5074> A_IWL<5073> A_IWL<5072> A_IWL<5071> A_IWL<5070> A_IWL<5069> A_IWL<5068> A_IWL<5067> A_IWL<5066> A_IWL<5065> A_IWL<5064> A_IWL<5063> A_IWL<5062> A_IWL<5061> A_IWL<5060> A_IWL<5059> A_IWL<5058> A_IWL<5057> A_IWL<5056> A_IWL<5055> A_IWL<5054> A_IWL<5053> A_IWL<5052> A_IWL<5051> A_IWL<5050> A_IWL<5049> A_IWL<5048> A_IWL<5047> A_IWL<5046> A_IWL<5045> A_IWL<5044> A_IWL<5043> A_IWL<5042> A_IWL<5041> A_IWL<5040> A_IWL<5039> A_IWL<5038> A_IWL<5037> A_IWL<5036> A_IWL<5035> A_IWL<5034> A_IWL<5033> A_IWL<5032> A_IWL<5031> A_IWL<5030> A_IWL<5029> A_IWL<5028> A_IWL<5027> A_IWL<5026> A_IWL<5025> A_IWL<5024> A_IWL<5023> A_IWL<5022> A_IWL<5021> A_IWL<5020> A_IWL<5019> A_IWL<5018> A_IWL<5017> A_IWL<5016> A_IWL<5015> A_IWL<5014> A_IWL<5013> A_IWL<5012> A_IWL<5011> A_IWL<5010> A_IWL<5009> A_IWL<5008> A_IWL<5007> A_IWL<5006> A_IWL<5005> A_IWL<5004> A_IWL<5003> A_IWL<5002> A_IWL<5001> A_IWL<5000> A_IWL<4999> A_IWL<4998> A_IWL<4997> A_IWL<4996> A_IWL<4995> A_IWL<4994> A_IWL<4993> A_IWL<4992> A_IWL<4991> A_IWL<4990> A_IWL<4989> A_IWL<4988> A_IWL<4987> A_IWL<4986> A_IWL<4985> A_IWL<4984> A_IWL<4983> A_IWL<4982> A_IWL<4981> A_IWL<4980> A_IWL<4979> A_IWL<4978> A_IWL<4977> A_IWL<4976> A_IWL<4975> A_IWL<4974> A_IWL<4973> A_IWL<4972> A_IWL<4971> A_IWL<4970> A_IWL<4969> A_IWL<4968> A_IWL<4967> A_IWL<4966> A_IWL<4965> A_IWL<4964> A_IWL<4963> A_IWL<4962> A_IWL<4961> A_IWL<4960> A_IWL<4959> A_IWL<4958> A_IWL<4957> A_IWL<4956> A_IWL<4955> A_IWL<4954> A_IWL<4953> A_IWL<4952> A_IWL<4951> A_IWL<4950> A_IWL<4949> A_IWL<4948> A_IWL<4947> A_IWL<4946> A_IWL<4945> A_IWL<4944> A_IWL<4943> A_IWL<4942> A_IWL<4941> A_IWL<4940> A_IWL<4939> A_IWL<4938> A_IWL<4937> A_IWL<4936> A_IWL<4935> A_IWL<4934> A_IWL<4933> A_IWL<4932> A_IWL<4931> A_IWL<4930> A_IWL<4929> A_IWL<4928> A_IWL<4927> A_IWL<4926> A_IWL<4925> A_IWL<4924> A_IWL<4923> A_IWL<4922> A_IWL<4921> A_IWL<4920> A_IWL<4919> A_IWL<4918> A_IWL<4917> A_IWL<4916> A_IWL<4915> A_IWL<4914> A_IWL<4913> A_IWL<4912> A_IWL<4911> A_IWL<4910> A_IWL<4909> A_IWL<4908> A_IWL<4907> A_IWL<4906> A_IWL<4905> A_IWL<4904> A_IWL<4903> A_IWL<4902> A_IWL<4901> A_IWL<4900> A_IWL<4899> A_IWL<4898> A_IWL<4897> A_IWL<4896> A_IWL<4895> A_IWL<4894> A_IWL<4893> A_IWL<4892> A_IWL<4891> A_IWL<4890> A_IWL<4889> A_IWL<4888> A_IWL<4887> A_IWL<4886> A_IWL<4885> A_IWL<4884> A_IWL<4883> A_IWL<4882> A_IWL<4881> A_IWL<4880> A_IWL<4879> A_IWL<4878> A_IWL<4877> A_IWL<4876> A_IWL<4875> A_IWL<4874> A_IWL<4873> A_IWL<4872> A_IWL<4871> A_IWL<4870> A_IWL<4869> A_IWL<4868> A_IWL<4867> A_IWL<4866> A_IWL<4865> A_IWL<4864> A_IWL<4863> A_IWL<4862> A_IWL<4861> A_IWL<4860> A_IWL<4859> A_IWL<4858> A_IWL<4857> A_IWL<4856> A_IWL<4855> A_IWL<4854> A_IWL<4853> A_IWL<4852> A_IWL<4851> A_IWL<4850> A_IWL<4849> A_IWL<4848> A_IWL<4847> A_IWL<4846> A_IWL<4845> A_IWL<4844> A_IWL<4843> A_IWL<4842> A_IWL<4841> A_IWL<4840> A_IWL<4839> A_IWL<4838> A_IWL<4837> A_IWL<4836> A_IWL<4835> A_IWL<4834> A_IWL<4833> A_IWL<4832> A_IWL<4831> A_IWL<4830> A_IWL<4829> A_IWL<4828> A_IWL<4827> A_IWL<4826> A_IWL<4825> A_IWL<4824> A_IWL<4823> A_IWL<4822> A_IWL<4821> A_IWL<4820> A_IWL<4819> A_IWL<4818> A_IWL<4817> A_IWL<4816> A_IWL<4815> A_IWL<4814> A_IWL<4813> A_IWL<4812> A_IWL<4811> A_IWL<4810> A_IWL<4809> A_IWL<4808> A_IWL<4807> A_IWL<4806> A_IWL<4805> A_IWL<4804> A_IWL<4803> A_IWL<4802> A_IWL<4801> A_IWL<4800> A_IWL<4799> A_IWL<4798> A_IWL<4797> A_IWL<4796> A_IWL<4795> A_IWL<4794> A_IWL<4793> A_IWL<4792> A_IWL<4791> A_IWL<4790> A_IWL<4789> A_IWL<4788> A_IWL<4787> A_IWL<4786> A_IWL<4785> A_IWL<4784> A_IWL<4783> A_IWL<4782> A_IWL<4781> A_IWL<4780> A_IWL<4779> A_IWL<4778> A_IWL<4777> A_IWL<4776> A_IWL<4775> A_IWL<4774> A_IWL<4773> A_IWL<4772> A_IWL<4771> A_IWL<4770> A_IWL<4769> A_IWL<4768> A_IWL<4767> A_IWL<4766> A_IWL<4765> A_IWL<4764> A_IWL<4763> A_IWL<4762> A_IWL<4761> A_IWL<4760> A_IWL<4759> A_IWL<4758> A_IWL<4757> A_IWL<4756> A_IWL<4755> A_IWL<4754> A_IWL<4753> A_IWL<4752> A_IWL<4751> A_IWL<4750> A_IWL<4749> A_IWL<4748> A_IWL<4747> A_IWL<4746> A_IWL<4745> A_IWL<4744> A_IWL<4743> A_IWL<4742> A_IWL<4741> A_IWL<4740> A_IWL<4739> A_IWL<4738> A_IWL<4737> A_IWL<4736> A_IWL<4735> A_IWL<4734> A_IWL<4733> A_IWL<4732> A_IWL<4731> A_IWL<4730> A_IWL<4729> A_IWL<4728> A_IWL<4727> A_IWL<4726> A_IWL<4725> A_IWL<4724> A_IWL<4723> A_IWL<4722> A_IWL<4721> A_IWL<4720> A_IWL<4719> A_IWL<4718> A_IWL<4717> A_IWL<4716> A_IWL<4715> A_IWL<4714> A_IWL<4713> A_IWL<4712> A_IWL<4711> A_IWL<4710> A_IWL<4709> A_IWL<4708> A_IWL<4707> A_IWL<4706> A_IWL<4705> A_IWL<4704> A_IWL<4703> A_IWL<4702> A_IWL<4701> A_IWL<4700> A_IWL<4699> A_IWL<4698> A_IWL<4697> A_IWL<4696> A_IWL<4695> A_IWL<4694> A_IWL<4693> A_IWL<4692> A_IWL<4691> A_IWL<4690> A_IWL<4689> A_IWL<4688> A_IWL<4687> A_IWL<4686> A_IWL<4685> A_IWL<4684> A_IWL<4683> A_IWL<4682> A_IWL<4681> A_IWL<4680> A_IWL<4679> A_IWL<4678> A_IWL<4677> A_IWL<4676> A_IWL<4675> A_IWL<4674> A_IWL<4673> A_IWL<4672> A_IWL<4671> A_IWL<4670> A_IWL<4669> A_IWL<4668> A_IWL<4667> A_IWL<4666> A_IWL<4665> A_IWL<4664> A_IWL<4663> A_IWL<4662> A_IWL<4661> A_IWL<4660> A_IWL<4659> A_IWL<4658> A_IWL<4657> A_IWL<4656> A_IWL<4655> A_IWL<4654> A_IWL<4653> A_IWL<4652> A_IWL<4651> A_IWL<4650> A_IWL<4649> A_IWL<4648> A_IWL<4647> A_IWL<4646> A_IWL<4645> A_IWL<4644> A_IWL<4643> A_IWL<4642> A_IWL<4641> A_IWL<4640> A_IWL<4639> A_IWL<4638> A_IWL<4637> A_IWL<4636> A_IWL<4635> A_IWL<4634> A_IWL<4633> A_IWL<4632> A_IWL<4631> A_IWL<4630> A_IWL<4629> A_IWL<4628> A_IWL<4627> A_IWL<4626> A_IWL<4625> A_IWL<4624> A_IWL<4623> A_IWL<4622> A_IWL<4621> A_IWL<4620> A_IWL<4619> A_IWL<4618> A_IWL<4617> A_IWL<4616> A_IWL<4615> A_IWL<4614> A_IWL<4613> A_IWL<4612> A_IWL<4611> A_IWL<4610> A_IWL<4609> A_IWL<4608> A_IWL<5631> A_IWL<5630> A_IWL<5629> A_IWL<5628> A_IWL<5627> A_IWL<5626> A_IWL<5625> A_IWL<5624> A_IWL<5623> A_IWL<5622> A_IWL<5621> A_IWL<5620> A_IWL<5619> A_IWL<5618> A_IWL<5617> A_IWL<5616> A_IWL<5615> A_IWL<5614> A_IWL<5613> A_IWL<5612> A_IWL<5611> A_IWL<5610> A_IWL<5609> A_IWL<5608> A_IWL<5607> A_IWL<5606> A_IWL<5605> A_IWL<5604> A_IWL<5603> A_IWL<5602> A_IWL<5601> A_IWL<5600> A_IWL<5599> A_IWL<5598> A_IWL<5597> A_IWL<5596> A_IWL<5595> A_IWL<5594> A_IWL<5593> A_IWL<5592> A_IWL<5591> A_IWL<5590> A_IWL<5589> A_IWL<5588> A_IWL<5587> A_IWL<5586> A_IWL<5585> A_IWL<5584> A_IWL<5583> A_IWL<5582> A_IWL<5581> A_IWL<5580> A_IWL<5579> A_IWL<5578> A_IWL<5577> A_IWL<5576> A_IWL<5575> A_IWL<5574> A_IWL<5573> A_IWL<5572> A_IWL<5571> A_IWL<5570> A_IWL<5569> A_IWL<5568> A_IWL<5567> A_IWL<5566> A_IWL<5565> A_IWL<5564> A_IWL<5563> A_IWL<5562> A_IWL<5561> A_IWL<5560> A_IWL<5559> A_IWL<5558> A_IWL<5557> A_IWL<5556> A_IWL<5555> A_IWL<5554> A_IWL<5553> A_IWL<5552> A_IWL<5551> A_IWL<5550> A_IWL<5549> A_IWL<5548> A_IWL<5547> A_IWL<5546> A_IWL<5545> A_IWL<5544> A_IWL<5543> A_IWL<5542> A_IWL<5541> A_IWL<5540> A_IWL<5539> A_IWL<5538> A_IWL<5537> A_IWL<5536> A_IWL<5535> A_IWL<5534> A_IWL<5533> A_IWL<5532> A_IWL<5531> A_IWL<5530> A_IWL<5529> A_IWL<5528> A_IWL<5527> A_IWL<5526> A_IWL<5525> A_IWL<5524> A_IWL<5523> A_IWL<5522> A_IWL<5521> A_IWL<5520> A_IWL<5519> A_IWL<5518> A_IWL<5517> A_IWL<5516> A_IWL<5515> A_IWL<5514> A_IWL<5513> A_IWL<5512> A_IWL<5511> A_IWL<5510> A_IWL<5509> A_IWL<5508> A_IWL<5507> A_IWL<5506> A_IWL<5505> A_IWL<5504> A_IWL<5503> A_IWL<5502> A_IWL<5501> A_IWL<5500> A_IWL<5499> A_IWL<5498> A_IWL<5497> A_IWL<5496> A_IWL<5495> A_IWL<5494> A_IWL<5493> A_IWL<5492> A_IWL<5491> A_IWL<5490> A_IWL<5489> A_IWL<5488> A_IWL<5487> A_IWL<5486> A_IWL<5485> A_IWL<5484> A_IWL<5483> A_IWL<5482> A_IWL<5481> A_IWL<5480> A_IWL<5479> A_IWL<5478> A_IWL<5477> A_IWL<5476> A_IWL<5475> A_IWL<5474> A_IWL<5473> A_IWL<5472> A_IWL<5471> A_IWL<5470> A_IWL<5469> A_IWL<5468> A_IWL<5467> A_IWL<5466> A_IWL<5465> A_IWL<5464> A_IWL<5463> A_IWL<5462> A_IWL<5461> A_IWL<5460> A_IWL<5459> A_IWL<5458> A_IWL<5457> A_IWL<5456> A_IWL<5455> A_IWL<5454> A_IWL<5453> A_IWL<5452> A_IWL<5451> A_IWL<5450> A_IWL<5449> A_IWL<5448> A_IWL<5447> A_IWL<5446> A_IWL<5445> A_IWL<5444> A_IWL<5443> A_IWL<5442> A_IWL<5441> A_IWL<5440> A_IWL<5439> A_IWL<5438> A_IWL<5437> A_IWL<5436> A_IWL<5435> A_IWL<5434> A_IWL<5433> A_IWL<5432> A_IWL<5431> A_IWL<5430> A_IWL<5429> A_IWL<5428> A_IWL<5427> A_IWL<5426> A_IWL<5425> A_IWL<5424> A_IWL<5423> A_IWL<5422> A_IWL<5421> A_IWL<5420> A_IWL<5419> A_IWL<5418> A_IWL<5417> A_IWL<5416> A_IWL<5415> A_IWL<5414> A_IWL<5413> A_IWL<5412> A_IWL<5411> A_IWL<5410> A_IWL<5409> A_IWL<5408> A_IWL<5407> A_IWL<5406> A_IWL<5405> A_IWL<5404> A_IWL<5403> A_IWL<5402> A_IWL<5401> A_IWL<5400> A_IWL<5399> A_IWL<5398> A_IWL<5397> A_IWL<5396> A_IWL<5395> A_IWL<5394> A_IWL<5393> A_IWL<5392> A_IWL<5391> A_IWL<5390> A_IWL<5389> A_IWL<5388> A_IWL<5387> A_IWL<5386> A_IWL<5385> A_IWL<5384> A_IWL<5383> A_IWL<5382> A_IWL<5381> A_IWL<5380> A_IWL<5379> A_IWL<5378> A_IWL<5377> A_IWL<5376> A_IWL<5375> A_IWL<5374> A_IWL<5373> A_IWL<5372> A_IWL<5371> A_IWL<5370> A_IWL<5369> A_IWL<5368> A_IWL<5367> A_IWL<5366> A_IWL<5365> A_IWL<5364> A_IWL<5363> A_IWL<5362> A_IWL<5361> A_IWL<5360> A_IWL<5359> A_IWL<5358> A_IWL<5357> A_IWL<5356> A_IWL<5355> A_IWL<5354> A_IWL<5353> A_IWL<5352> A_IWL<5351> A_IWL<5350> A_IWL<5349> A_IWL<5348> A_IWL<5347> A_IWL<5346> A_IWL<5345> A_IWL<5344> A_IWL<5343> A_IWL<5342> A_IWL<5341> A_IWL<5340> A_IWL<5339> A_IWL<5338> A_IWL<5337> A_IWL<5336> A_IWL<5335> A_IWL<5334> A_IWL<5333> A_IWL<5332> A_IWL<5331> A_IWL<5330> A_IWL<5329> A_IWL<5328> A_IWL<5327> A_IWL<5326> A_IWL<5325> A_IWL<5324> A_IWL<5323> A_IWL<5322> A_IWL<5321> A_IWL<5320> A_IWL<5319> A_IWL<5318> A_IWL<5317> A_IWL<5316> A_IWL<5315> A_IWL<5314> A_IWL<5313> A_IWL<5312> A_IWL<5311> A_IWL<5310> A_IWL<5309> A_IWL<5308> A_IWL<5307> A_IWL<5306> A_IWL<5305> A_IWL<5304> A_IWL<5303> A_IWL<5302> A_IWL<5301> A_IWL<5300> A_IWL<5299> A_IWL<5298> A_IWL<5297> A_IWL<5296> A_IWL<5295> A_IWL<5294> A_IWL<5293> A_IWL<5292> A_IWL<5291> A_IWL<5290> A_IWL<5289> A_IWL<5288> A_IWL<5287> A_IWL<5286> A_IWL<5285> A_IWL<5284> A_IWL<5283> A_IWL<5282> A_IWL<5281> A_IWL<5280> A_IWL<5279> A_IWL<5278> A_IWL<5277> A_IWL<5276> A_IWL<5275> A_IWL<5274> A_IWL<5273> A_IWL<5272> A_IWL<5271> A_IWL<5270> A_IWL<5269> A_IWL<5268> A_IWL<5267> A_IWL<5266> A_IWL<5265> A_IWL<5264> A_IWL<5263> A_IWL<5262> A_IWL<5261> A_IWL<5260> A_IWL<5259> A_IWL<5258> A_IWL<5257> A_IWL<5256> A_IWL<5255> A_IWL<5254> A_IWL<5253> A_IWL<5252> A_IWL<5251> A_IWL<5250> A_IWL<5249> A_IWL<5248> A_IWL<5247> A_IWL<5246> A_IWL<5245> A_IWL<5244> A_IWL<5243> A_IWL<5242> A_IWL<5241> A_IWL<5240> A_IWL<5239> A_IWL<5238> A_IWL<5237> A_IWL<5236> A_IWL<5235> A_IWL<5234> A_IWL<5233> A_IWL<5232> A_IWL<5231> A_IWL<5230> A_IWL<5229> A_IWL<5228> A_IWL<5227> A_IWL<5226> A_IWL<5225> A_IWL<5224> A_IWL<5223> A_IWL<5222> A_IWL<5221> A_IWL<5220> A_IWL<5219> A_IWL<5218> A_IWL<5217> A_IWL<5216> A_IWL<5215> A_IWL<5214> A_IWL<5213> A_IWL<5212> A_IWL<5211> A_IWL<5210> A_IWL<5209> A_IWL<5208> A_IWL<5207> A_IWL<5206> A_IWL<5205> A_IWL<5204> A_IWL<5203> A_IWL<5202> A_IWL<5201> A_IWL<5200> A_IWL<5199> A_IWL<5198> A_IWL<5197> A_IWL<5196> A_IWL<5195> A_IWL<5194> A_IWL<5193> A_IWL<5192> A_IWL<5191> A_IWL<5190> A_IWL<5189> A_IWL<5188> A_IWL<5187> A_IWL<5186> A_IWL<5185> A_IWL<5184> A_IWL<5183> A_IWL<5182> A_IWL<5181> A_IWL<5180> A_IWL<5179> A_IWL<5178> A_IWL<5177> A_IWL<5176> A_IWL<5175> A_IWL<5174> A_IWL<5173> A_IWL<5172> A_IWL<5171> A_IWL<5170> A_IWL<5169> A_IWL<5168> A_IWL<5167> A_IWL<5166> A_IWL<5165> A_IWL<5164> A_IWL<5163> A_IWL<5162> A_IWL<5161> A_IWL<5160> A_IWL<5159> A_IWL<5158> A_IWL<5157> A_IWL<5156> A_IWL<5155> A_IWL<5154> A_IWL<5153> A_IWL<5152> A_IWL<5151> A_IWL<5150> A_IWL<5149> A_IWL<5148> A_IWL<5147> A_IWL<5146> A_IWL<5145> A_IWL<5144> A_IWL<5143> A_IWL<5142> A_IWL<5141> A_IWL<5140> A_IWL<5139> A_IWL<5138> A_IWL<5137> A_IWL<5136> A_IWL<5135> A_IWL<5134> A_IWL<5133> A_IWL<5132> A_IWL<5131> A_IWL<5130> A_IWL<5129> A_IWL<5128> A_IWL<5127> A_IWL<5126> A_IWL<5125> A_IWL<5124> A_IWL<5123> A_IWL<5122> A_IWL<5121> A_IWL<5120> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<9> A_BLC<19> A_BLC<18> A_BLC_TOP<19> A_BLC_TOP<18> A_BLT<19> A_BLT<18> A_BLT_TOP<19> A_BLT_TOP<18> A_IWL<4607> A_IWL<4606> A_IWL<4605> A_IWL<4604> A_IWL<4603> A_IWL<4602> A_IWL<4601> A_IWL<4600> A_IWL<4599> A_IWL<4598> A_IWL<4597> A_IWL<4596> A_IWL<4595> A_IWL<4594> A_IWL<4593> A_IWL<4592> A_IWL<4591> A_IWL<4590> A_IWL<4589> A_IWL<4588> A_IWL<4587> A_IWL<4586> A_IWL<4585> A_IWL<4584> A_IWL<4583> A_IWL<4582> A_IWL<4581> A_IWL<4580> A_IWL<4579> A_IWL<4578> A_IWL<4577> A_IWL<4576> A_IWL<4575> A_IWL<4574> A_IWL<4573> A_IWL<4572> A_IWL<4571> A_IWL<4570> A_IWL<4569> A_IWL<4568> A_IWL<4567> A_IWL<4566> A_IWL<4565> A_IWL<4564> A_IWL<4563> A_IWL<4562> A_IWL<4561> A_IWL<4560> A_IWL<4559> A_IWL<4558> A_IWL<4557> A_IWL<4556> A_IWL<4555> A_IWL<4554> A_IWL<4553> A_IWL<4552> A_IWL<4551> A_IWL<4550> A_IWL<4549> A_IWL<4548> A_IWL<4547> A_IWL<4546> A_IWL<4545> A_IWL<4544> A_IWL<4543> A_IWL<4542> A_IWL<4541> A_IWL<4540> A_IWL<4539> A_IWL<4538> A_IWL<4537> A_IWL<4536> A_IWL<4535> A_IWL<4534> A_IWL<4533> A_IWL<4532> A_IWL<4531> A_IWL<4530> A_IWL<4529> A_IWL<4528> A_IWL<4527> A_IWL<4526> A_IWL<4525> A_IWL<4524> A_IWL<4523> A_IWL<4522> A_IWL<4521> A_IWL<4520> A_IWL<4519> A_IWL<4518> A_IWL<4517> A_IWL<4516> A_IWL<4515> A_IWL<4514> A_IWL<4513> A_IWL<4512> A_IWL<4511> A_IWL<4510> A_IWL<4509> A_IWL<4508> A_IWL<4507> A_IWL<4506> A_IWL<4505> A_IWL<4504> A_IWL<4503> A_IWL<4502> A_IWL<4501> A_IWL<4500> A_IWL<4499> A_IWL<4498> A_IWL<4497> A_IWL<4496> A_IWL<4495> A_IWL<4494> A_IWL<4493> A_IWL<4492> A_IWL<4491> A_IWL<4490> A_IWL<4489> A_IWL<4488> A_IWL<4487> A_IWL<4486> A_IWL<4485> A_IWL<4484> A_IWL<4483> A_IWL<4482> A_IWL<4481> A_IWL<4480> A_IWL<4479> A_IWL<4478> A_IWL<4477> A_IWL<4476> A_IWL<4475> A_IWL<4474> A_IWL<4473> A_IWL<4472> A_IWL<4471> A_IWL<4470> A_IWL<4469> A_IWL<4468> A_IWL<4467> A_IWL<4466> A_IWL<4465> A_IWL<4464> A_IWL<4463> A_IWL<4462> A_IWL<4461> A_IWL<4460> A_IWL<4459> A_IWL<4458> A_IWL<4457> A_IWL<4456> A_IWL<4455> A_IWL<4454> A_IWL<4453> A_IWL<4452> A_IWL<4451> A_IWL<4450> A_IWL<4449> A_IWL<4448> A_IWL<4447> A_IWL<4446> A_IWL<4445> A_IWL<4444> A_IWL<4443> A_IWL<4442> A_IWL<4441> A_IWL<4440> A_IWL<4439> A_IWL<4438> A_IWL<4437> A_IWL<4436> A_IWL<4435> A_IWL<4434> A_IWL<4433> A_IWL<4432> A_IWL<4431> A_IWL<4430> A_IWL<4429> A_IWL<4428> A_IWL<4427> A_IWL<4426> A_IWL<4425> A_IWL<4424> A_IWL<4423> A_IWL<4422> A_IWL<4421> A_IWL<4420> A_IWL<4419> A_IWL<4418> A_IWL<4417> A_IWL<4416> A_IWL<4415> A_IWL<4414> A_IWL<4413> A_IWL<4412> A_IWL<4411> A_IWL<4410> A_IWL<4409> A_IWL<4408> A_IWL<4407> A_IWL<4406> A_IWL<4405> A_IWL<4404> A_IWL<4403> A_IWL<4402> A_IWL<4401> A_IWL<4400> A_IWL<4399> A_IWL<4398> A_IWL<4397> A_IWL<4396> A_IWL<4395> A_IWL<4394> A_IWL<4393> A_IWL<4392> A_IWL<4391> A_IWL<4390> A_IWL<4389> A_IWL<4388> A_IWL<4387> A_IWL<4386> A_IWL<4385> A_IWL<4384> A_IWL<4383> A_IWL<4382> A_IWL<4381> A_IWL<4380> A_IWL<4379> A_IWL<4378> A_IWL<4377> A_IWL<4376> A_IWL<4375> A_IWL<4374> A_IWL<4373> A_IWL<4372> A_IWL<4371> A_IWL<4370> A_IWL<4369> A_IWL<4368> A_IWL<4367> A_IWL<4366> A_IWL<4365> A_IWL<4364> A_IWL<4363> A_IWL<4362> A_IWL<4361> A_IWL<4360> A_IWL<4359> A_IWL<4358> A_IWL<4357> A_IWL<4356> A_IWL<4355> A_IWL<4354> A_IWL<4353> A_IWL<4352> A_IWL<4351> A_IWL<4350> A_IWL<4349> A_IWL<4348> A_IWL<4347> A_IWL<4346> A_IWL<4345> A_IWL<4344> A_IWL<4343> A_IWL<4342> A_IWL<4341> A_IWL<4340> A_IWL<4339> A_IWL<4338> A_IWL<4337> A_IWL<4336> A_IWL<4335> A_IWL<4334> A_IWL<4333> A_IWL<4332> A_IWL<4331> A_IWL<4330> A_IWL<4329> A_IWL<4328> A_IWL<4327> A_IWL<4326> A_IWL<4325> A_IWL<4324> A_IWL<4323> A_IWL<4322> A_IWL<4321> A_IWL<4320> A_IWL<4319> A_IWL<4318> A_IWL<4317> A_IWL<4316> A_IWL<4315> A_IWL<4314> A_IWL<4313> A_IWL<4312> A_IWL<4311> A_IWL<4310> A_IWL<4309> A_IWL<4308> A_IWL<4307> A_IWL<4306> A_IWL<4305> A_IWL<4304> A_IWL<4303> A_IWL<4302> A_IWL<4301> A_IWL<4300> A_IWL<4299> A_IWL<4298> A_IWL<4297> A_IWL<4296> A_IWL<4295> A_IWL<4294> A_IWL<4293> A_IWL<4292> A_IWL<4291> A_IWL<4290> A_IWL<4289> A_IWL<4288> A_IWL<4287> A_IWL<4286> A_IWL<4285> A_IWL<4284> A_IWL<4283> A_IWL<4282> A_IWL<4281> A_IWL<4280> A_IWL<4279> A_IWL<4278> A_IWL<4277> A_IWL<4276> A_IWL<4275> A_IWL<4274> A_IWL<4273> A_IWL<4272> A_IWL<4271> A_IWL<4270> A_IWL<4269> A_IWL<4268> A_IWL<4267> A_IWL<4266> A_IWL<4265> A_IWL<4264> A_IWL<4263> A_IWL<4262> A_IWL<4261> A_IWL<4260> A_IWL<4259> A_IWL<4258> A_IWL<4257> A_IWL<4256> A_IWL<4255> A_IWL<4254> A_IWL<4253> A_IWL<4252> A_IWL<4251> A_IWL<4250> A_IWL<4249> A_IWL<4248> A_IWL<4247> A_IWL<4246> A_IWL<4245> A_IWL<4244> A_IWL<4243> A_IWL<4242> A_IWL<4241> A_IWL<4240> A_IWL<4239> A_IWL<4238> A_IWL<4237> A_IWL<4236> A_IWL<4235> A_IWL<4234> A_IWL<4233> A_IWL<4232> A_IWL<4231> A_IWL<4230> A_IWL<4229> A_IWL<4228> A_IWL<4227> A_IWL<4226> A_IWL<4225> A_IWL<4224> A_IWL<4223> A_IWL<4222> A_IWL<4221> A_IWL<4220> A_IWL<4219> A_IWL<4218> A_IWL<4217> A_IWL<4216> A_IWL<4215> A_IWL<4214> A_IWL<4213> A_IWL<4212> A_IWL<4211> A_IWL<4210> A_IWL<4209> A_IWL<4208> A_IWL<4207> A_IWL<4206> A_IWL<4205> A_IWL<4204> A_IWL<4203> A_IWL<4202> A_IWL<4201> A_IWL<4200> A_IWL<4199> A_IWL<4198> A_IWL<4197> A_IWL<4196> A_IWL<4195> A_IWL<4194> A_IWL<4193> A_IWL<4192> A_IWL<4191> A_IWL<4190> A_IWL<4189> A_IWL<4188> A_IWL<4187> A_IWL<4186> A_IWL<4185> A_IWL<4184> A_IWL<4183> A_IWL<4182> A_IWL<4181> A_IWL<4180> A_IWL<4179> A_IWL<4178> A_IWL<4177> A_IWL<4176> A_IWL<4175> A_IWL<4174> A_IWL<4173> A_IWL<4172> A_IWL<4171> A_IWL<4170> A_IWL<4169> A_IWL<4168> A_IWL<4167> A_IWL<4166> A_IWL<4165> A_IWL<4164> A_IWL<4163> A_IWL<4162> A_IWL<4161> A_IWL<4160> A_IWL<4159> A_IWL<4158> A_IWL<4157> A_IWL<4156> A_IWL<4155> A_IWL<4154> A_IWL<4153> A_IWL<4152> A_IWL<4151> A_IWL<4150> A_IWL<4149> A_IWL<4148> A_IWL<4147> A_IWL<4146> A_IWL<4145> A_IWL<4144> A_IWL<4143> A_IWL<4142> A_IWL<4141> A_IWL<4140> A_IWL<4139> A_IWL<4138> A_IWL<4137> A_IWL<4136> A_IWL<4135> A_IWL<4134> A_IWL<4133> A_IWL<4132> A_IWL<4131> A_IWL<4130> A_IWL<4129> A_IWL<4128> A_IWL<4127> A_IWL<4126> A_IWL<4125> A_IWL<4124> A_IWL<4123> A_IWL<4122> A_IWL<4121> A_IWL<4120> A_IWL<4119> A_IWL<4118> A_IWL<4117> A_IWL<4116> A_IWL<4115> A_IWL<4114> A_IWL<4113> A_IWL<4112> A_IWL<4111> A_IWL<4110> A_IWL<4109> A_IWL<4108> A_IWL<4107> A_IWL<4106> A_IWL<4105> A_IWL<4104> A_IWL<4103> A_IWL<4102> A_IWL<4101> A_IWL<4100> A_IWL<4099> A_IWL<4098> A_IWL<4097> A_IWL<4096> A_IWL<5119> A_IWL<5118> A_IWL<5117> A_IWL<5116> A_IWL<5115> A_IWL<5114> A_IWL<5113> A_IWL<5112> A_IWL<5111> A_IWL<5110> A_IWL<5109> A_IWL<5108> A_IWL<5107> A_IWL<5106> A_IWL<5105> A_IWL<5104> A_IWL<5103> A_IWL<5102> A_IWL<5101> A_IWL<5100> A_IWL<5099> A_IWL<5098> A_IWL<5097> A_IWL<5096> A_IWL<5095> A_IWL<5094> A_IWL<5093> A_IWL<5092> A_IWL<5091> A_IWL<5090> A_IWL<5089> A_IWL<5088> A_IWL<5087> A_IWL<5086> A_IWL<5085> A_IWL<5084> A_IWL<5083> A_IWL<5082> A_IWL<5081> A_IWL<5080> A_IWL<5079> A_IWL<5078> A_IWL<5077> A_IWL<5076> A_IWL<5075> A_IWL<5074> A_IWL<5073> A_IWL<5072> A_IWL<5071> A_IWL<5070> A_IWL<5069> A_IWL<5068> A_IWL<5067> A_IWL<5066> A_IWL<5065> A_IWL<5064> A_IWL<5063> A_IWL<5062> A_IWL<5061> A_IWL<5060> A_IWL<5059> A_IWL<5058> A_IWL<5057> A_IWL<5056> A_IWL<5055> A_IWL<5054> A_IWL<5053> A_IWL<5052> A_IWL<5051> A_IWL<5050> A_IWL<5049> A_IWL<5048> A_IWL<5047> A_IWL<5046> A_IWL<5045> A_IWL<5044> A_IWL<5043> A_IWL<5042> A_IWL<5041> A_IWL<5040> A_IWL<5039> A_IWL<5038> A_IWL<5037> A_IWL<5036> A_IWL<5035> A_IWL<5034> A_IWL<5033> A_IWL<5032> A_IWL<5031> A_IWL<5030> A_IWL<5029> A_IWL<5028> A_IWL<5027> A_IWL<5026> A_IWL<5025> A_IWL<5024> A_IWL<5023> A_IWL<5022> A_IWL<5021> A_IWL<5020> A_IWL<5019> A_IWL<5018> A_IWL<5017> A_IWL<5016> A_IWL<5015> A_IWL<5014> A_IWL<5013> A_IWL<5012> A_IWL<5011> A_IWL<5010> A_IWL<5009> A_IWL<5008> A_IWL<5007> A_IWL<5006> A_IWL<5005> A_IWL<5004> A_IWL<5003> A_IWL<5002> A_IWL<5001> A_IWL<5000> A_IWL<4999> A_IWL<4998> A_IWL<4997> A_IWL<4996> A_IWL<4995> A_IWL<4994> A_IWL<4993> A_IWL<4992> A_IWL<4991> A_IWL<4990> A_IWL<4989> A_IWL<4988> A_IWL<4987> A_IWL<4986> A_IWL<4985> A_IWL<4984> A_IWL<4983> A_IWL<4982> A_IWL<4981> A_IWL<4980> A_IWL<4979> A_IWL<4978> A_IWL<4977> A_IWL<4976> A_IWL<4975> A_IWL<4974> A_IWL<4973> A_IWL<4972> A_IWL<4971> A_IWL<4970> A_IWL<4969> A_IWL<4968> A_IWL<4967> A_IWL<4966> A_IWL<4965> A_IWL<4964> A_IWL<4963> A_IWL<4962> A_IWL<4961> A_IWL<4960> A_IWL<4959> A_IWL<4958> A_IWL<4957> A_IWL<4956> A_IWL<4955> A_IWL<4954> A_IWL<4953> A_IWL<4952> A_IWL<4951> A_IWL<4950> A_IWL<4949> A_IWL<4948> A_IWL<4947> A_IWL<4946> A_IWL<4945> A_IWL<4944> A_IWL<4943> A_IWL<4942> A_IWL<4941> A_IWL<4940> A_IWL<4939> A_IWL<4938> A_IWL<4937> A_IWL<4936> A_IWL<4935> A_IWL<4934> A_IWL<4933> A_IWL<4932> A_IWL<4931> A_IWL<4930> A_IWL<4929> A_IWL<4928> A_IWL<4927> A_IWL<4926> A_IWL<4925> A_IWL<4924> A_IWL<4923> A_IWL<4922> A_IWL<4921> A_IWL<4920> A_IWL<4919> A_IWL<4918> A_IWL<4917> A_IWL<4916> A_IWL<4915> A_IWL<4914> A_IWL<4913> A_IWL<4912> A_IWL<4911> A_IWL<4910> A_IWL<4909> A_IWL<4908> A_IWL<4907> A_IWL<4906> A_IWL<4905> A_IWL<4904> A_IWL<4903> A_IWL<4902> A_IWL<4901> A_IWL<4900> A_IWL<4899> A_IWL<4898> A_IWL<4897> A_IWL<4896> A_IWL<4895> A_IWL<4894> A_IWL<4893> A_IWL<4892> A_IWL<4891> A_IWL<4890> A_IWL<4889> A_IWL<4888> A_IWL<4887> A_IWL<4886> A_IWL<4885> A_IWL<4884> A_IWL<4883> A_IWL<4882> A_IWL<4881> A_IWL<4880> A_IWL<4879> A_IWL<4878> A_IWL<4877> A_IWL<4876> A_IWL<4875> A_IWL<4874> A_IWL<4873> A_IWL<4872> A_IWL<4871> A_IWL<4870> A_IWL<4869> A_IWL<4868> A_IWL<4867> A_IWL<4866> A_IWL<4865> A_IWL<4864> A_IWL<4863> A_IWL<4862> A_IWL<4861> A_IWL<4860> A_IWL<4859> A_IWL<4858> A_IWL<4857> A_IWL<4856> A_IWL<4855> A_IWL<4854> A_IWL<4853> A_IWL<4852> A_IWL<4851> A_IWL<4850> A_IWL<4849> A_IWL<4848> A_IWL<4847> A_IWL<4846> A_IWL<4845> A_IWL<4844> A_IWL<4843> A_IWL<4842> A_IWL<4841> A_IWL<4840> A_IWL<4839> A_IWL<4838> A_IWL<4837> A_IWL<4836> A_IWL<4835> A_IWL<4834> A_IWL<4833> A_IWL<4832> A_IWL<4831> A_IWL<4830> A_IWL<4829> A_IWL<4828> A_IWL<4827> A_IWL<4826> A_IWL<4825> A_IWL<4824> A_IWL<4823> A_IWL<4822> A_IWL<4821> A_IWL<4820> A_IWL<4819> A_IWL<4818> A_IWL<4817> A_IWL<4816> A_IWL<4815> A_IWL<4814> A_IWL<4813> A_IWL<4812> A_IWL<4811> A_IWL<4810> A_IWL<4809> A_IWL<4808> A_IWL<4807> A_IWL<4806> A_IWL<4805> A_IWL<4804> A_IWL<4803> A_IWL<4802> A_IWL<4801> A_IWL<4800> A_IWL<4799> A_IWL<4798> A_IWL<4797> A_IWL<4796> A_IWL<4795> A_IWL<4794> A_IWL<4793> A_IWL<4792> A_IWL<4791> A_IWL<4790> A_IWL<4789> A_IWL<4788> A_IWL<4787> A_IWL<4786> A_IWL<4785> A_IWL<4784> A_IWL<4783> A_IWL<4782> A_IWL<4781> A_IWL<4780> A_IWL<4779> A_IWL<4778> A_IWL<4777> A_IWL<4776> A_IWL<4775> A_IWL<4774> A_IWL<4773> A_IWL<4772> A_IWL<4771> A_IWL<4770> A_IWL<4769> A_IWL<4768> A_IWL<4767> A_IWL<4766> A_IWL<4765> A_IWL<4764> A_IWL<4763> A_IWL<4762> A_IWL<4761> A_IWL<4760> A_IWL<4759> A_IWL<4758> A_IWL<4757> A_IWL<4756> A_IWL<4755> A_IWL<4754> A_IWL<4753> A_IWL<4752> A_IWL<4751> A_IWL<4750> A_IWL<4749> A_IWL<4748> A_IWL<4747> A_IWL<4746> A_IWL<4745> A_IWL<4744> A_IWL<4743> A_IWL<4742> A_IWL<4741> A_IWL<4740> A_IWL<4739> A_IWL<4738> A_IWL<4737> A_IWL<4736> A_IWL<4735> A_IWL<4734> A_IWL<4733> A_IWL<4732> A_IWL<4731> A_IWL<4730> A_IWL<4729> A_IWL<4728> A_IWL<4727> A_IWL<4726> A_IWL<4725> A_IWL<4724> A_IWL<4723> A_IWL<4722> A_IWL<4721> A_IWL<4720> A_IWL<4719> A_IWL<4718> A_IWL<4717> A_IWL<4716> A_IWL<4715> A_IWL<4714> A_IWL<4713> A_IWL<4712> A_IWL<4711> A_IWL<4710> A_IWL<4709> A_IWL<4708> A_IWL<4707> A_IWL<4706> A_IWL<4705> A_IWL<4704> A_IWL<4703> A_IWL<4702> A_IWL<4701> A_IWL<4700> A_IWL<4699> A_IWL<4698> A_IWL<4697> A_IWL<4696> A_IWL<4695> A_IWL<4694> A_IWL<4693> A_IWL<4692> A_IWL<4691> A_IWL<4690> A_IWL<4689> A_IWL<4688> A_IWL<4687> A_IWL<4686> A_IWL<4685> A_IWL<4684> A_IWL<4683> A_IWL<4682> A_IWL<4681> A_IWL<4680> A_IWL<4679> A_IWL<4678> A_IWL<4677> A_IWL<4676> A_IWL<4675> A_IWL<4674> A_IWL<4673> A_IWL<4672> A_IWL<4671> A_IWL<4670> A_IWL<4669> A_IWL<4668> A_IWL<4667> A_IWL<4666> A_IWL<4665> A_IWL<4664> A_IWL<4663> A_IWL<4662> A_IWL<4661> A_IWL<4660> A_IWL<4659> A_IWL<4658> A_IWL<4657> A_IWL<4656> A_IWL<4655> A_IWL<4654> A_IWL<4653> A_IWL<4652> A_IWL<4651> A_IWL<4650> A_IWL<4649> A_IWL<4648> A_IWL<4647> A_IWL<4646> A_IWL<4645> A_IWL<4644> A_IWL<4643> A_IWL<4642> A_IWL<4641> A_IWL<4640> A_IWL<4639> A_IWL<4638> A_IWL<4637> A_IWL<4636> A_IWL<4635> A_IWL<4634> A_IWL<4633> A_IWL<4632> A_IWL<4631> A_IWL<4630> A_IWL<4629> A_IWL<4628> A_IWL<4627> A_IWL<4626> A_IWL<4625> A_IWL<4624> A_IWL<4623> A_IWL<4622> A_IWL<4621> A_IWL<4620> A_IWL<4619> A_IWL<4618> A_IWL<4617> A_IWL<4616> A_IWL<4615> A_IWL<4614> A_IWL<4613> A_IWL<4612> A_IWL<4611> A_IWL<4610> A_IWL<4609> A_IWL<4608> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<8> A_BLC<17> A_BLC<16> A_BLC_TOP<17> A_BLC_TOP<16> A_BLT<17> A_BLT<16> A_BLT_TOP<17> A_BLT_TOP<16> A_IWL<4095> A_IWL<4094> A_IWL<4093> A_IWL<4092> A_IWL<4091> A_IWL<4090> A_IWL<4089> A_IWL<4088> A_IWL<4087> A_IWL<4086> A_IWL<4085> A_IWL<4084> A_IWL<4083> A_IWL<4082> A_IWL<4081> A_IWL<4080> A_IWL<4079> A_IWL<4078> A_IWL<4077> A_IWL<4076> A_IWL<4075> A_IWL<4074> A_IWL<4073> A_IWL<4072> A_IWL<4071> A_IWL<4070> A_IWL<4069> A_IWL<4068> A_IWL<4067> A_IWL<4066> A_IWL<4065> A_IWL<4064> A_IWL<4063> A_IWL<4062> A_IWL<4061> A_IWL<4060> A_IWL<4059> A_IWL<4058> A_IWL<4057> A_IWL<4056> A_IWL<4055> A_IWL<4054> A_IWL<4053> A_IWL<4052> A_IWL<4051> A_IWL<4050> A_IWL<4049> A_IWL<4048> A_IWL<4047> A_IWL<4046> A_IWL<4045> A_IWL<4044> A_IWL<4043> A_IWL<4042> A_IWL<4041> A_IWL<4040> A_IWL<4039> A_IWL<4038> A_IWL<4037> A_IWL<4036> A_IWL<4035> A_IWL<4034> A_IWL<4033> A_IWL<4032> A_IWL<4031> A_IWL<4030> A_IWL<4029> A_IWL<4028> A_IWL<4027> A_IWL<4026> A_IWL<4025> A_IWL<4024> A_IWL<4023> A_IWL<4022> A_IWL<4021> A_IWL<4020> A_IWL<4019> A_IWL<4018> A_IWL<4017> A_IWL<4016> A_IWL<4015> A_IWL<4014> A_IWL<4013> A_IWL<4012> A_IWL<4011> A_IWL<4010> A_IWL<4009> A_IWL<4008> A_IWL<4007> A_IWL<4006> A_IWL<4005> A_IWL<4004> A_IWL<4003> A_IWL<4002> A_IWL<4001> A_IWL<4000> A_IWL<3999> A_IWL<3998> A_IWL<3997> A_IWL<3996> A_IWL<3995> A_IWL<3994> A_IWL<3993> A_IWL<3992> A_IWL<3991> A_IWL<3990> A_IWL<3989> A_IWL<3988> A_IWL<3987> A_IWL<3986> A_IWL<3985> A_IWL<3984> A_IWL<3983> A_IWL<3982> A_IWL<3981> A_IWL<3980> A_IWL<3979> A_IWL<3978> A_IWL<3977> A_IWL<3976> A_IWL<3975> A_IWL<3974> A_IWL<3973> A_IWL<3972> A_IWL<3971> A_IWL<3970> A_IWL<3969> A_IWL<3968> A_IWL<3967> A_IWL<3966> A_IWL<3965> A_IWL<3964> A_IWL<3963> A_IWL<3962> A_IWL<3961> A_IWL<3960> A_IWL<3959> A_IWL<3958> A_IWL<3957> A_IWL<3956> A_IWL<3955> A_IWL<3954> A_IWL<3953> A_IWL<3952> A_IWL<3951> A_IWL<3950> A_IWL<3949> A_IWL<3948> A_IWL<3947> A_IWL<3946> A_IWL<3945> A_IWL<3944> A_IWL<3943> A_IWL<3942> A_IWL<3941> A_IWL<3940> A_IWL<3939> A_IWL<3938> A_IWL<3937> A_IWL<3936> A_IWL<3935> A_IWL<3934> A_IWL<3933> A_IWL<3932> A_IWL<3931> A_IWL<3930> A_IWL<3929> A_IWL<3928> A_IWL<3927> A_IWL<3926> A_IWL<3925> A_IWL<3924> A_IWL<3923> A_IWL<3922> A_IWL<3921> A_IWL<3920> A_IWL<3919> A_IWL<3918> A_IWL<3917> A_IWL<3916> A_IWL<3915> A_IWL<3914> A_IWL<3913> A_IWL<3912> A_IWL<3911> A_IWL<3910> A_IWL<3909> A_IWL<3908> A_IWL<3907> A_IWL<3906> A_IWL<3905> A_IWL<3904> A_IWL<3903> A_IWL<3902> A_IWL<3901> A_IWL<3900> A_IWL<3899> A_IWL<3898> A_IWL<3897> A_IWL<3896> A_IWL<3895> A_IWL<3894> A_IWL<3893> A_IWL<3892> A_IWL<3891> A_IWL<3890> A_IWL<3889> A_IWL<3888> A_IWL<3887> A_IWL<3886> A_IWL<3885> A_IWL<3884> A_IWL<3883> A_IWL<3882> A_IWL<3881> A_IWL<3880> A_IWL<3879> A_IWL<3878> A_IWL<3877> A_IWL<3876> A_IWL<3875> A_IWL<3874> A_IWL<3873> A_IWL<3872> A_IWL<3871> A_IWL<3870> A_IWL<3869> A_IWL<3868> A_IWL<3867> A_IWL<3866> A_IWL<3865> A_IWL<3864> A_IWL<3863> A_IWL<3862> A_IWL<3861> A_IWL<3860> A_IWL<3859> A_IWL<3858> A_IWL<3857> A_IWL<3856> A_IWL<3855> A_IWL<3854> A_IWL<3853> A_IWL<3852> A_IWL<3851> A_IWL<3850> A_IWL<3849> A_IWL<3848> A_IWL<3847> A_IWL<3846> A_IWL<3845> A_IWL<3844> A_IWL<3843> A_IWL<3842> A_IWL<3841> A_IWL<3840> A_IWL<3839> A_IWL<3838> A_IWL<3837> A_IWL<3836> A_IWL<3835> A_IWL<3834> A_IWL<3833> A_IWL<3832> A_IWL<3831> A_IWL<3830> A_IWL<3829> A_IWL<3828> A_IWL<3827> A_IWL<3826> A_IWL<3825> A_IWL<3824> A_IWL<3823> A_IWL<3822> A_IWL<3821> A_IWL<3820> A_IWL<3819> A_IWL<3818> A_IWL<3817> A_IWL<3816> A_IWL<3815> A_IWL<3814> A_IWL<3813> A_IWL<3812> A_IWL<3811> A_IWL<3810> A_IWL<3809> A_IWL<3808> A_IWL<3807> A_IWL<3806> A_IWL<3805> A_IWL<3804> A_IWL<3803> A_IWL<3802> A_IWL<3801> A_IWL<3800> A_IWL<3799> A_IWL<3798> A_IWL<3797> A_IWL<3796> A_IWL<3795> A_IWL<3794> A_IWL<3793> A_IWL<3792> A_IWL<3791> A_IWL<3790> A_IWL<3789> A_IWL<3788> A_IWL<3787> A_IWL<3786> A_IWL<3785> A_IWL<3784> A_IWL<3783> A_IWL<3782> A_IWL<3781> A_IWL<3780> A_IWL<3779> A_IWL<3778> A_IWL<3777> A_IWL<3776> A_IWL<3775> A_IWL<3774> A_IWL<3773> A_IWL<3772> A_IWL<3771> A_IWL<3770> A_IWL<3769> A_IWL<3768> A_IWL<3767> A_IWL<3766> A_IWL<3765> A_IWL<3764> A_IWL<3763> A_IWL<3762> A_IWL<3761> A_IWL<3760> A_IWL<3759> A_IWL<3758> A_IWL<3757> A_IWL<3756> A_IWL<3755> A_IWL<3754> A_IWL<3753> A_IWL<3752> A_IWL<3751> A_IWL<3750> A_IWL<3749> A_IWL<3748> A_IWL<3747> A_IWL<3746> A_IWL<3745> A_IWL<3744> A_IWL<3743> A_IWL<3742> A_IWL<3741> A_IWL<3740> A_IWL<3739> A_IWL<3738> A_IWL<3737> A_IWL<3736> A_IWL<3735> A_IWL<3734> A_IWL<3733> A_IWL<3732> A_IWL<3731> A_IWL<3730> A_IWL<3729> A_IWL<3728> A_IWL<3727> A_IWL<3726> A_IWL<3725> A_IWL<3724> A_IWL<3723> A_IWL<3722> A_IWL<3721> A_IWL<3720> A_IWL<3719> A_IWL<3718> A_IWL<3717> A_IWL<3716> A_IWL<3715> A_IWL<3714> A_IWL<3713> A_IWL<3712> A_IWL<3711> A_IWL<3710> A_IWL<3709> A_IWL<3708> A_IWL<3707> A_IWL<3706> A_IWL<3705> A_IWL<3704> A_IWL<3703> A_IWL<3702> A_IWL<3701> A_IWL<3700> A_IWL<3699> A_IWL<3698> A_IWL<3697> A_IWL<3696> A_IWL<3695> A_IWL<3694> A_IWL<3693> A_IWL<3692> A_IWL<3691> A_IWL<3690> A_IWL<3689> A_IWL<3688> A_IWL<3687> A_IWL<3686> A_IWL<3685> A_IWL<3684> A_IWL<3683> A_IWL<3682> A_IWL<3681> A_IWL<3680> A_IWL<3679> A_IWL<3678> A_IWL<3677> A_IWL<3676> A_IWL<3675> A_IWL<3674> A_IWL<3673> A_IWL<3672> A_IWL<3671> A_IWL<3670> A_IWL<3669> A_IWL<3668> A_IWL<3667> A_IWL<3666> A_IWL<3665> A_IWL<3664> A_IWL<3663> A_IWL<3662> A_IWL<3661> A_IWL<3660> A_IWL<3659> A_IWL<3658> A_IWL<3657> A_IWL<3656> A_IWL<3655> A_IWL<3654> A_IWL<3653> A_IWL<3652> A_IWL<3651> A_IWL<3650> A_IWL<3649> A_IWL<3648> A_IWL<3647> A_IWL<3646> A_IWL<3645> A_IWL<3644> A_IWL<3643> A_IWL<3642> A_IWL<3641> A_IWL<3640> A_IWL<3639> A_IWL<3638> A_IWL<3637> A_IWL<3636> A_IWL<3635> A_IWL<3634> A_IWL<3633> A_IWL<3632> A_IWL<3631> A_IWL<3630> A_IWL<3629> A_IWL<3628> A_IWL<3627> A_IWL<3626> A_IWL<3625> A_IWL<3624> A_IWL<3623> A_IWL<3622> A_IWL<3621> A_IWL<3620> A_IWL<3619> A_IWL<3618> A_IWL<3617> A_IWL<3616> A_IWL<3615> A_IWL<3614> A_IWL<3613> A_IWL<3612> A_IWL<3611> A_IWL<3610> A_IWL<3609> A_IWL<3608> A_IWL<3607> A_IWL<3606> A_IWL<3605> A_IWL<3604> A_IWL<3603> A_IWL<3602> A_IWL<3601> A_IWL<3600> A_IWL<3599> A_IWL<3598> A_IWL<3597> A_IWL<3596> A_IWL<3595> A_IWL<3594> A_IWL<3593> A_IWL<3592> A_IWL<3591> A_IWL<3590> A_IWL<3589> A_IWL<3588> A_IWL<3587> A_IWL<3586> A_IWL<3585> A_IWL<3584> A_IWL<4607> A_IWL<4606> A_IWL<4605> A_IWL<4604> A_IWL<4603> A_IWL<4602> A_IWL<4601> A_IWL<4600> A_IWL<4599> A_IWL<4598> A_IWL<4597> A_IWL<4596> A_IWL<4595> A_IWL<4594> A_IWL<4593> A_IWL<4592> A_IWL<4591> A_IWL<4590> A_IWL<4589> A_IWL<4588> A_IWL<4587> A_IWL<4586> A_IWL<4585> A_IWL<4584> A_IWL<4583> A_IWL<4582> A_IWL<4581> A_IWL<4580> A_IWL<4579> A_IWL<4578> A_IWL<4577> A_IWL<4576> A_IWL<4575> A_IWL<4574> A_IWL<4573> A_IWL<4572> A_IWL<4571> A_IWL<4570> A_IWL<4569> A_IWL<4568> A_IWL<4567> A_IWL<4566> A_IWL<4565> A_IWL<4564> A_IWL<4563> A_IWL<4562> A_IWL<4561> A_IWL<4560> A_IWL<4559> A_IWL<4558> A_IWL<4557> A_IWL<4556> A_IWL<4555> A_IWL<4554> A_IWL<4553> A_IWL<4552> A_IWL<4551> A_IWL<4550> A_IWL<4549> A_IWL<4548> A_IWL<4547> A_IWL<4546> A_IWL<4545> A_IWL<4544> A_IWL<4543> A_IWL<4542> A_IWL<4541> A_IWL<4540> A_IWL<4539> A_IWL<4538> A_IWL<4537> A_IWL<4536> A_IWL<4535> A_IWL<4534> A_IWL<4533> A_IWL<4532> A_IWL<4531> A_IWL<4530> A_IWL<4529> A_IWL<4528> A_IWL<4527> A_IWL<4526> A_IWL<4525> A_IWL<4524> A_IWL<4523> A_IWL<4522> A_IWL<4521> A_IWL<4520> A_IWL<4519> A_IWL<4518> A_IWL<4517> A_IWL<4516> A_IWL<4515> A_IWL<4514> A_IWL<4513> A_IWL<4512> A_IWL<4511> A_IWL<4510> A_IWL<4509> A_IWL<4508> A_IWL<4507> A_IWL<4506> A_IWL<4505> A_IWL<4504> A_IWL<4503> A_IWL<4502> A_IWL<4501> A_IWL<4500> A_IWL<4499> A_IWL<4498> A_IWL<4497> A_IWL<4496> A_IWL<4495> A_IWL<4494> A_IWL<4493> A_IWL<4492> A_IWL<4491> A_IWL<4490> A_IWL<4489> A_IWL<4488> A_IWL<4487> A_IWL<4486> A_IWL<4485> A_IWL<4484> A_IWL<4483> A_IWL<4482> A_IWL<4481> A_IWL<4480> A_IWL<4479> A_IWL<4478> A_IWL<4477> A_IWL<4476> A_IWL<4475> A_IWL<4474> A_IWL<4473> A_IWL<4472> A_IWL<4471> A_IWL<4470> A_IWL<4469> A_IWL<4468> A_IWL<4467> A_IWL<4466> A_IWL<4465> A_IWL<4464> A_IWL<4463> A_IWL<4462> A_IWL<4461> A_IWL<4460> A_IWL<4459> A_IWL<4458> A_IWL<4457> A_IWL<4456> A_IWL<4455> A_IWL<4454> A_IWL<4453> A_IWL<4452> A_IWL<4451> A_IWL<4450> A_IWL<4449> A_IWL<4448> A_IWL<4447> A_IWL<4446> A_IWL<4445> A_IWL<4444> A_IWL<4443> A_IWL<4442> A_IWL<4441> A_IWL<4440> A_IWL<4439> A_IWL<4438> A_IWL<4437> A_IWL<4436> A_IWL<4435> A_IWL<4434> A_IWL<4433> A_IWL<4432> A_IWL<4431> A_IWL<4430> A_IWL<4429> A_IWL<4428> A_IWL<4427> A_IWL<4426> A_IWL<4425> A_IWL<4424> A_IWL<4423> A_IWL<4422> A_IWL<4421> A_IWL<4420> A_IWL<4419> A_IWL<4418> A_IWL<4417> A_IWL<4416> A_IWL<4415> A_IWL<4414> A_IWL<4413> A_IWL<4412> A_IWL<4411> A_IWL<4410> A_IWL<4409> A_IWL<4408> A_IWL<4407> A_IWL<4406> A_IWL<4405> A_IWL<4404> A_IWL<4403> A_IWL<4402> A_IWL<4401> A_IWL<4400> A_IWL<4399> A_IWL<4398> A_IWL<4397> A_IWL<4396> A_IWL<4395> A_IWL<4394> A_IWL<4393> A_IWL<4392> A_IWL<4391> A_IWL<4390> A_IWL<4389> A_IWL<4388> A_IWL<4387> A_IWL<4386> A_IWL<4385> A_IWL<4384> A_IWL<4383> A_IWL<4382> A_IWL<4381> A_IWL<4380> A_IWL<4379> A_IWL<4378> A_IWL<4377> A_IWL<4376> A_IWL<4375> A_IWL<4374> A_IWL<4373> A_IWL<4372> A_IWL<4371> A_IWL<4370> A_IWL<4369> A_IWL<4368> A_IWL<4367> A_IWL<4366> A_IWL<4365> A_IWL<4364> A_IWL<4363> A_IWL<4362> A_IWL<4361> A_IWL<4360> A_IWL<4359> A_IWL<4358> A_IWL<4357> A_IWL<4356> A_IWL<4355> A_IWL<4354> A_IWL<4353> A_IWL<4352> A_IWL<4351> A_IWL<4350> A_IWL<4349> A_IWL<4348> A_IWL<4347> A_IWL<4346> A_IWL<4345> A_IWL<4344> A_IWL<4343> A_IWL<4342> A_IWL<4341> A_IWL<4340> A_IWL<4339> A_IWL<4338> A_IWL<4337> A_IWL<4336> A_IWL<4335> A_IWL<4334> A_IWL<4333> A_IWL<4332> A_IWL<4331> A_IWL<4330> A_IWL<4329> A_IWL<4328> A_IWL<4327> A_IWL<4326> A_IWL<4325> A_IWL<4324> A_IWL<4323> A_IWL<4322> A_IWL<4321> A_IWL<4320> A_IWL<4319> A_IWL<4318> A_IWL<4317> A_IWL<4316> A_IWL<4315> A_IWL<4314> A_IWL<4313> A_IWL<4312> A_IWL<4311> A_IWL<4310> A_IWL<4309> A_IWL<4308> A_IWL<4307> A_IWL<4306> A_IWL<4305> A_IWL<4304> A_IWL<4303> A_IWL<4302> A_IWL<4301> A_IWL<4300> A_IWL<4299> A_IWL<4298> A_IWL<4297> A_IWL<4296> A_IWL<4295> A_IWL<4294> A_IWL<4293> A_IWL<4292> A_IWL<4291> A_IWL<4290> A_IWL<4289> A_IWL<4288> A_IWL<4287> A_IWL<4286> A_IWL<4285> A_IWL<4284> A_IWL<4283> A_IWL<4282> A_IWL<4281> A_IWL<4280> A_IWL<4279> A_IWL<4278> A_IWL<4277> A_IWL<4276> A_IWL<4275> A_IWL<4274> A_IWL<4273> A_IWL<4272> A_IWL<4271> A_IWL<4270> A_IWL<4269> A_IWL<4268> A_IWL<4267> A_IWL<4266> A_IWL<4265> A_IWL<4264> A_IWL<4263> A_IWL<4262> A_IWL<4261> A_IWL<4260> A_IWL<4259> A_IWL<4258> A_IWL<4257> A_IWL<4256> A_IWL<4255> A_IWL<4254> A_IWL<4253> A_IWL<4252> A_IWL<4251> A_IWL<4250> A_IWL<4249> A_IWL<4248> A_IWL<4247> A_IWL<4246> A_IWL<4245> A_IWL<4244> A_IWL<4243> A_IWL<4242> A_IWL<4241> A_IWL<4240> A_IWL<4239> A_IWL<4238> A_IWL<4237> A_IWL<4236> A_IWL<4235> A_IWL<4234> A_IWL<4233> A_IWL<4232> A_IWL<4231> A_IWL<4230> A_IWL<4229> A_IWL<4228> A_IWL<4227> A_IWL<4226> A_IWL<4225> A_IWL<4224> A_IWL<4223> A_IWL<4222> A_IWL<4221> A_IWL<4220> A_IWL<4219> A_IWL<4218> A_IWL<4217> A_IWL<4216> A_IWL<4215> A_IWL<4214> A_IWL<4213> A_IWL<4212> A_IWL<4211> A_IWL<4210> A_IWL<4209> A_IWL<4208> A_IWL<4207> A_IWL<4206> A_IWL<4205> A_IWL<4204> A_IWL<4203> A_IWL<4202> A_IWL<4201> A_IWL<4200> A_IWL<4199> A_IWL<4198> A_IWL<4197> A_IWL<4196> A_IWL<4195> A_IWL<4194> A_IWL<4193> A_IWL<4192> A_IWL<4191> A_IWL<4190> A_IWL<4189> A_IWL<4188> A_IWL<4187> A_IWL<4186> A_IWL<4185> A_IWL<4184> A_IWL<4183> A_IWL<4182> A_IWL<4181> A_IWL<4180> A_IWL<4179> A_IWL<4178> A_IWL<4177> A_IWL<4176> A_IWL<4175> A_IWL<4174> A_IWL<4173> A_IWL<4172> A_IWL<4171> A_IWL<4170> A_IWL<4169> A_IWL<4168> A_IWL<4167> A_IWL<4166> A_IWL<4165> A_IWL<4164> A_IWL<4163> A_IWL<4162> A_IWL<4161> A_IWL<4160> A_IWL<4159> A_IWL<4158> A_IWL<4157> A_IWL<4156> A_IWL<4155> A_IWL<4154> A_IWL<4153> A_IWL<4152> A_IWL<4151> A_IWL<4150> A_IWL<4149> A_IWL<4148> A_IWL<4147> A_IWL<4146> A_IWL<4145> A_IWL<4144> A_IWL<4143> A_IWL<4142> A_IWL<4141> A_IWL<4140> A_IWL<4139> A_IWL<4138> A_IWL<4137> A_IWL<4136> A_IWL<4135> A_IWL<4134> A_IWL<4133> A_IWL<4132> A_IWL<4131> A_IWL<4130> A_IWL<4129> A_IWL<4128> A_IWL<4127> A_IWL<4126> A_IWL<4125> A_IWL<4124> A_IWL<4123> A_IWL<4122> A_IWL<4121> A_IWL<4120> A_IWL<4119> A_IWL<4118> A_IWL<4117> A_IWL<4116> A_IWL<4115> A_IWL<4114> A_IWL<4113> A_IWL<4112> A_IWL<4111> A_IWL<4110> A_IWL<4109> A_IWL<4108> A_IWL<4107> A_IWL<4106> A_IWL<4105> A_IWL<4104> A_IWL<4103> A_IWL<4102> A_IWL<4101> A_IWL<4100> A_IWL<4099> A_IWL<4098> A_IWL<4097> A_IWL<4096> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<7> A_BLC<15> A_BLC<14> A_BLC_TOP<15> A_BLC_TOP<14> A_BLT<15> A_BLT<14> A_BLT_TOP<15> A_BLT_TOP<14> A_IWL<3583> A_IWL<3582> A_IWL<3581> A_IWL<3580> A_IWL<3579> A_IWL<3578> A_IWL<3577> A_IWL<3576> A_IWL<3575> A_IWL<3574> A_IWL<3573> A_IWL<3572> A_IWL<3571> A_IWL<3570> A_IWL<3569> A_IWL<3568> A_IWL<3567> A_IWL<3566> A_IWL<3565> A_IWL<3564> A_IWL<3563> A_IWL<3562> A_IWL<3561> A_IWL<3560> A_IWL<3559> A_IWL<3558> A_IWL<3557> A_IWL<3556> A_IWL<3555> A_IWL<3554> A_IWL<3553> A_IWL<3552> A_IWL<3551> A_IWL<3550> A_IWL<3549> A_IWL<3548> A_IWL<3547> A_IWL<3546> A_IWL<3545> A_IWL<3544> A_IWL<3543> A_IWL<3542> A_IWL<3541> A_IWL<3540> A_IWL<3539> A_IWL<3538> A_IWL<3537> A_IWL<3536> A_IWL<3535> A_IWL<3534> A_IWL<3533> A_IWL<3532> A_IWL<3531> A_IWL<3530> A_IWL<3529> A_IWL<3528> A_IWL<3527> A_IWL<3526> A_IWL<3525> A_IWL<3524> A_IWL<3523> A_IWL<3522> A_IWL<3521> A_IWL<3520> A_IWL<3519> A_IWL<3518> A_IWL<3517> A_IWL<3516> A_IWL<3515> A_IWL<3514> A_IWL<3513> A_IWL<3512> A_IWL<3511> A_IWL<3510> A_IWL<3509> A_IWL<3508> A_IWL<3507> A_IWL<3506> A_IWL<3505> A_IWL<3504> A_IWL<3503> A_IWL<3502> A_IWL<3501> A_IWL<3500> A_IWL<3499> A_IWL<3498> A_IWL<3497> A_IWL<3496> A_IWL<3495> A_IWL<3494> A_IWL<3493> A_IWL<3492> A_IWL<3491> A_IWL<3490> A_IWL<3489> A_IWL<3488> A_IWL<3487> A_IWL<3486> A_IWL<3485> A_IWL<3484> A_IWL<3483> A_IWL<3482> A_IWL<3481> A_IWL<3480> A_IWL<3479> A_IWL<3478> A_IWL<3477> A_IWL<3476> A_IWL<3475> A_IWL<3474> A_IWL<3473> A_IWL<3472> A_IWL<3471> A_IWL<3470> A_IWL<3469> A_IWL<3468> A_IWL<3467> A_IWL<3466> A_IWL<3465> A_IWL<3464> A_IWL<3463> A_IWL<3462> A_IWL<3461> A_IWL<3460> A_IWL<3459> A_IWL<3458> A_IWL<3457> A_IWL<3456> A_IWL<3455> A_IWL<3454> A_IWL<3453> A_IWL<3452> A_IWL<3451> A_IWL<3450> A_IWL<3449> A_IWL<3448> A_IWL<3447> A_IWL<3446> A_IWL<3445> A_IWL<3444> A_IWL<3443> A_IWL<3442> A_IWL<3441> A_IWL<3440> A_IWL<3439> A_IWL<3438> A_IWL<3437> A_IWL<3436> A_IWL<3435> A_IWL<3434> A_IWL<3433> A_IWL<3432> A_IWL<3431> A_IWL<3430> A_IWL<3429> A_IWL<3428> A_IWL<3427> A_IWL<3426> A_IWL<3425> A_IWL<3424> A_IWL<3423> A_IWL<3422> A_IWL<3421> A_IWL<3420> A_IWL<3419> A_IWL<3418> A_IWL<3417> A_IWL<3416> A_IWL<3415> A_IWL<3414> A_IWL<3413> A_IWL<3412> A_IWL<3411> A_IWL<3410> A_IWL<3409> A_IWL<3408> A_IWL<3407> A_IWL<3406> A_IWL<3405> A_IWL<3404> A_IWL<3403> A_IWL<3402> A_IWL<3401> A_IWL<3400> A_IWL<3399> A_IWL<3398> A_IWL<3397> A_IWL<3396> A_IWL<3395> A_IWL<3394> A_IWL<3393> A_IWL<3392> A_IWL<3391> A_IWL<3390> A_IWL<3389> A_IWL<3388> A_IWL<3387> A_IWL<3386> A_IWL<3385> A_IWL<3384> A_IWL<3383> A_IWL<3382> A_IWL<3381> A_IWL<3380> A_IWL<3379> A_IWL<3378> A_IWL<3377> A_IWL<3376> A_IWL<3375> A_IWL<3374> A_IWL<3373> A_IWL<3372> A_IWL<3371> A_IWL<3370> A_IWL<3369> A_IWL<3368> A_IWL<3367> A_IWL<3366> A_IWL<3365> A_IWL<3364> A_IWL<3363> A_IWL<3362> A_IWL<3361> A_IWL<3360> A_IWL<3359> A_IWL<3358> A_IWL<3357> A_IWL<3356> A_IWL<3355> A_IWL<3354> A_IWL<3353> A_IWL<3352> A_IWL<3351> A_IWL<3350> A_IWL<3349> A_IWL<3348> A_IWL<3347> A_IWL<3346> A_IWL<3345> A_IWL<3344> A_IWL<3343> A_IWL<3342> A_IWL<3341> A_IWL<3340> A_IWL<3339> A_IWL<3338> A_IWL<3337> A_IWL<3336> A_IWL<3335> A_IWL<3334> A_IWL<3333> A_IWL<3332> A_IWL<3331> A_IWL<3330> A_IWL<3329> A_IWL<3328> A_IWL<3327> A_IWL<3326> A_IWL<3325> A_IWL<3324> A_IWL<3323> A_IWL<3322> A_IWL<3321> A_IWL<3320> A_IWL<3319> A_IWL<3318> A_IWL<3317> A_IWL<3316> A_IWL<3315> A_IWL<3314> A_IWL<3313> A_IWL<3312> A_IWL<3311> A_IWL<3310> A_IWL<3309> A_IWL<3308> A_IWL<3307> A_IWL<3306> A_IWL<3305> A_IWL<3304> A_IWL<3303> A_IWL<3302> A_IWL<3301> A_IWL<3300> A_IWL<3299> A_IWL<3298> A_IWL<3297> A_IWL<3296> A_IWL<3295> A_IWL<3294> A_IWL<3293> A_IWL<3292> A_IWL<3291> A_IWL<3290> A_IWL<3289> A_IWL<3288> A_IWL<3287> A_IWL<3286> A_IWL<3285> A_IWL<3284> A_IWL<3283> A_IWL<3282> A_IWL<3281> A_IWL<3280> A_IWL<3279> A_IWL<3278> A_IWL<3277> A_IWL<3276> A_IWL<3275> A_IWL<3274> A_IWL<3273> A_IWL<3272> A_IWL<3271> A_IWL<3270> A_IWL<3269> A_IWL<3268> A_IWL<3267> A_IWL<3266> A_IWL<3265> A_IWL<3264> A_IWL<3263> A_IWL<3262> A_IWL<3261> A_IWL<3260> A_IWL<3259> A_IWL<3258> A_IWL<3257> A_IWL<3256> A_IWL<3255> A_IWL<3254> A_IWL<3253> A_IWL<3252> A_IWL<3251> A_IWL<3250> A_IWL<3249> A_IWL<3248> A_IWL<3247> A_IWL<3246> A_IWL<3245> A_IWL<3244> A_IWL<3243> A_IWL<3242> A_IWL<3241> A_IWL<3240> A_IWL<3239> A_IWL<3238> A_IWL<3237> A_IWL<3236> A_IWL<3235> A_IWL<3234> A_IWL<3233> A_IWL<3232> A_IWL<3231> A_IWL<3230> A_IWL<3229> A_IWL<3228> A_IWL<3227> A_IWL<3226> A_IWL<3225> A_IWL<3224> A_IWL<3223> A_IWL<3222> A_IWL<3221> A_IWL<3220> A_IWL<3219> A_IWL<3218> A_IWL<3217> A_IWL<3216> A_IWL<3215> A_IWL<3214> A_IWL<3213> A_IWL<3212> A_IWL<3211> A_IWL<3210> A_IWL<3209> A_IWL<3208> A_IWL<3207> A_IWL<3206> A_IWL<3205> A_IWL<3204> A_IWL<3203> A_IWL<3202> A_IWL<3201> A_IWL<3200> A_IWL<3199> A_IWL<3198> A_IWL<3197> A_IWL<3196> A_IWL<3195> A_IWL<3194> A_IWL<3193> A_IWL<3192> A_IWL<3191> A_IWL<3190> A_IWL<3189> A_IWL<3188> A_IWL<3187> A_IWL<3186> A_IWL<3185> A_IWL<3184> A_IWL<3183> A_IWL<3182> A_IWL<3181> A_IWL<3180> A_IWL<3179> A_IWL<3178> A_IWL<3177> A_IWL<3176> A_IWL<3175> A_IWL<3174> A_IWL<3173> A_IWL<3172> A_IWL<3171> A_IWL<3170> A_IWL<3169> A_IWL<3168> A_IWL<3167> A_IWL<3166> A_IWL<3165> A_IWL<3164> A_IWL<3163> A_IWL<3162> A_IWL<3161> A_IWL<3160> A_IWL<3159> A_IWL<3158> A_IWL<3157> A_IWL<3156> A_IWL<3155> A_IWL<3154> A_IWL<3153> A_IWL<3152> A_IWL<3151> A_IWL<3150> A_IWL<3149> A_IWL<3148> A_IWL<3147> A_IWL<3146> A_IWL<3145> A_IWL<3144> A_IWL<3143> A_IWL<3142> A_IWL<3141> A_IWL<3140> A_IWL<3139> A_IWL<3138> A_IWL<3137> A_IWL<3136> A_IWL<3135> A_IWL<3134> A_IWL<3133> A_IWL<3132> A_IWL<3131> A_IWL<3130> A_IWL<3129> A_IWL<3128> A_IWL<3127> A_IWL<3126> A_IWL<3125> A_IWL<3124> A_IWL<3123> A_IWL<3122> A_IWL<3121> A_IWL<3120> A_IWL<3119> A_IWL<3118> A_IWL<3117> A_IWL<3116> A_IWL<3115> A_IWL<3114> A_IWL<3113> A_IWL<3112> A_IWL<3111> A_IWL<3110> A_IWL<3109> A_IWL<3108> A_IWL<3107> A_IWL<3106> A_IWL<3105> A_IWL<3104> A_IWL<3103> A_IWL<3102> A_IWL<3101> A_IWL<3100> A_IWL<3099> A_IWL<3098> A_IWL<3097> A_IWL<3096> A_IWL<3095> A_IWL<3094> A_IWL<3093> A_IWL<3092> A_IWL<3091> A_IWL<3090> A_IWL<3089> A_IWL<3088> A_IWL<3087> A_IWL<3086> A_IWL<3085> A_IWL<3084> A_IWL<3083> A_IWL<3082> A_IWL<3081> A_IWL<3080> A_IWL<3079> A_IWL<3078> A_IWL<3077> A_IWL<3076> A_IWL<3075> A_IWL<3074> A_IWL<3073> A_IWL<3072> A_IWL<4095> A_IWL<4094> A_IWL<4093> A_IWL<4092> A_IWL<4091> A_IWL<4090> A_IWL<4089> A_IWL<4088> A_IWL<4087> A_IWL<4086> A_IWL<4085> A_IWL<4084> A_IWL<4083> A_IWL<4082> A_IWL<4081> A_IWL<4080> A_IWL<4079> A_IWL<4078> A_IWL<4077> A_IWL<4076> A_IWL<4075> A_IWL<4074> A_IWL<4073> A_IWL<4072> A_IWL<4071> A_IWL<4070> A_IWL<4069> A_IWL<4068> A_IWL<4067> A_IWL<4066> A_IWL<4065> A_IWL<4064> A_IWL<4063> A_IWL<4062> A_IWL<4061> A_IWL<4060> A_IWL<4059> A_IWL<4058> A_IWL<4057> A_IWL<4056> A_IWL<4055> A_IWL<4054> A_IWL<4053> A_IWL<4052> A_IWL<4051> A_IWL<4050> A_IWL<4049> A_IWL<4048> A_IWL<4047> A_IWL<4046> A_IWL<4045> A_IWL<4044> A_IWL<4043> A_IWL<4042> A_IWL<4041> A_IWL<4040> A_IWL<4039> A_IWL<4038> A_IWL<4037> A_IWL<4036> A_IWL<4035> A_IWL<4034> A_IWL<4033> A_IWL<4032> A_IWL<4031> A_IWL<4030> A_IWL<4029> A_IWL<4028> A_IWL<4027> A_IWL<4026> A_IWL<4025> A_IWL<4024> A_IWL<4023> A_IWL<4022> A_IWL<4021> A_IWL<4020> A_IWL<4019> A_IWL<4018> A_IWL<4017> A_IWL<4016> A_IWL<4015> A_IWL<4014> A_IWL<4013> A_IWL<4012> A_IWL<4011> A_IWL<4010> A_IWL<4009> A_IWL<4008> A_IWL<4007> A_IWL<4006> A_IWL<4005> A_IWL<4004> A_IWL<4003> A_IWL<4002> A_IWL<4001> A_IWL<4000> A_IWL<3999> A_IWL<3998> A_IWL<3997> A_IWL<3996> A_IWL<3995> A_IWL<3994> A_IWL<3993> A_IWL<3992> A_IWL<3991> A_IWL<3990> A_IWL<3989> A_IWL<3988> A_IWL<3987> A_IWL<3986> A_IWL<3985> A_IWL<3984> A_IWL<3983> A_IWL<3982> A_IWL<3981> A_IWL<3980> A_IWL<3979> A_IWL<3978> A_IWL<3977> A_IWL<3976> A_IWL<3975> A_IWL<3974> A_IWL<3973> A_IWL<3972> A_IWL<3971> A_IWL<3970> A_IWL<3969> A_IWL<3968> A_IWL<3967> A_IWL<3966> A_IWL<3965> A_IWL<3964> A_IWL<3963> A_IWL<3962> A_IWL<3961> A_IWL<3960> A_IWL<3959> A_IWL<3958> A_IWL<3957> A_IWL<3956> A_IWL<3955> A_IWL<3954> A_IWL<3953> A_IWL<3952> A_IWL<3951> A_IWL<3950> A_IWL<3949> A_IWL<3948> A_IWL<3947> A_IWL<3946> A_IWL<3945> A_IWL<3944> A_IWL<3943> A_IWL<3942> A_IWL<3941> A_IWL<3940> A_IWL<3939> A_IWL<3938> A_IWL<3937> A_IWL<3936> A_IWL<3935> A_IWL<3934> A_IWL<3933> A_IWL<3932> A_IWL<3931> A_IWL<3930> A_IWL<3929> A_IWL<3928> A_IWL<3927> A_IWL<3926> A_IWL<3925> A_IWL<3924> A_IWL<3923> A_IWL<3922> A_IWL<3921> A_IWL<3920> A_IWL<3919> A_IWL<3918> A_IWL<3917> A_IWL<3916> A_IWL<3915> A_IWL<3914> A_IWL<3913> A_IWL<3912> A_IWL<3911> A_IWL<3910> A_IWL<3909> A_IWL<3908> A_IWL<3907> A_IWL<3906> A_IWL<3905> A_IWL<3904> A_IWL<3903> A_IWL<3902> A_IWL<3901> A_IWL<3900> A_IWL<3899> A_IWL<3898> A_IWL<3897> A_IWL<3896> A_IWL<3895> A_IWL<3894> A_IWL<3893> A_IWL<3892> A_IWL<3891> A_IWL<3890> A_IWL<3889> A_IWL<3888> A_IWL<3887> A_IWL<3886> A_IWL<3885> A_IWL<3884> A_IWL<3883> A_IWL<3882> A_IWL<3881> A_IWL<3880> A_IWL<3879> A_IWL<3878> A_IWL<3877> A_IWL<3876> A_IWL<3875> A_IWL<3874> A_IWL<3873> A_IWL<3872> A_IWL<3871> A_IWL<3870> A_IWL<3869> A_IWL<3868> A_IWL<3867> A_IWL<3866> A_IWL<3865> A_IWL<3864> A_IWL<3863> A_IWL<3862> A_IWL<3861> A_IWL<3860> A_IWL<3859> A_IWL<3858> A_IWL<3857> A_IWL<3856> A_IWL<3855> A_IWL<3854> A_IWL<3853> A_IWL<3852> A_IWL<3851> A_IWL<3850> A_IWL<3849> A_IWL<3848> A_IWL<3847> A_IWL<3846> A_IWL<3845> A_IWL<3844> A_IWL<3843> A_IWL<3842> A_IWL<3841> A_IWL<3840> A_IWL<3839> A_IWL<3838> A_IWL<3837> A_IWL<3836> A_IWL<3835> A_IWL<3834> A_IWL<3833> A_IWL<3832> A_IWL<3831> A_IWL<3830> A_IWL<3829> A_IWL<3828> A_IWL<3827> A_IWL<3826> A_IWL<3825> A_IWL<3824> A_IWL<3823> A_IWL<3822> A_IWL<3821> A_IWL<3820> A_IWL<3819> A_IWL<3818> A_IWL<3817> A_IWL<3816> A_IWL<3815> A_IWL<3814> A_IWL<3813> A_IWL<3812> A_IWL<3811> A_IWL<3810> A_IWL<3809> A_IWL<3808> A_IWL<3807> A_IWL<3806> A_IWL<3805> A_IWL<3804> A_IWL<3803> A_IWL<3802> A_IWL<3801> A_IWL<3800> A_IWL<3799> A_IWL<3798> A_IWL<3797> A_IWL<3796> A_IWL<3795> A_IWL<3794> A_IWL<3793> A_IWL<3792> A_IWL<3791> A_IWL<3790> A_IWL<3789> A_IWL<3788> A_IWL<3787> A_IWL<3786> A_IWL<3785> A_IWL<3784> A_IWL<3783> A_IWL<3782> A_IWL<3781> A_IWL<3780> A_IWL<3779> A_IWL<3778> A_IWL<3777> A_IWL<3776> A_IWL<3775> A_IWL<3774> A_IWL<3773> A_IWL<3772> A_IWL<3771> A_IWL<3770> A_IWL<3769> A_IWL<3768> A_IWL<3767> A_IWL<3766> A_IWL<3765> A_IWL<3764> A_IWL<3763> A_IWL<3762> A_IWL<3761> A_IWL<3760> A_IWL<3759> A_IWL<3758> A_IWL<3757> A_IWL<3756> A_IWL<3755> A_IWL<3754> A_IWL<3753> A_IWL<3752> A_IWL<3751> A_IWL<3750> A_IWL<3749> A_IWL<3748> A_IWL<3747> A_IWL<3746> A_IWL<3745> A_IWL<3744> A_IWL<3743> A_IWL<3742> A_IWL<3741> A_IWL<3740> A_IWL<3739> A_IWL<3738> A_IWL<3737> A_IWL<3736> A_IWL<3735> A_IWL<3734> A_IWL<3733> A_IWL<3732> A_IWL<3731> A_IWL<3730> A_IWL<3729> A_IWL<3728> A_IWL<3727> A_IWL<3726> A_IWL<3725> A_IWL<3724> A_IWL<3723> A_IWL<3722> A_IWL<3721> A_IWL<3720> A_IWL<3719> A_IWL<3718> A_IWL<3717> A_IWL<3716> A_IWL<3715> A_IWL<3714> A_IWL<3713> A_IWL<3712> A_IWL<3711> A_IWL<3710> A_IWL<3709> A_IWL<3708> A_IWL<3707> A_IWL<3706> A_IWL<3705> A_IWL<3704> A_IWL<3703> A_IWL<3702> A_IWL<3701> A_IWL<3700> A_IWL<3699> A_IWL<3698> A_IWL<3697> A_IWL<3696> A_IWL<3695> A_IWL<3694> A_IWL<3693> A_IWL<3692> A_IWL<3691> A_IWL<3690> A_IWL<3689> A_IWL<3688> A_IWL<3687> A_IWL<3686> A_IWL<3685> A_IWL<3684> A_IWL<3683> A_IWL<3682> A_IWL<3681> A_IWL<3680> A_IWL<3679> A_IWL<3678> A_IWL<3677> A_IWL<3676> A_IWL<3675> A_IWL<3674> A_IWL<3673> A_IWL<3672> A_IWL<3671> A_IWL<3670> A_IWL<3669> A_IWL<3668> A_IWL<3667> A_IWL<3666> A_IWL<3665> A_IWL<3664> A_IWL<3663> A_IWL<3662> A_IWL<3661> A_IWL<3660> A_IWL<3659> A_IWL<3658> A_IWL<3657> A_IWL<3656> A_IWL<3655> A_IWL<3654> A_IWL<3653> A_IWL<3652> A_IWL<3651> A_IWL<3650> A_IWL<3649> A_IWL<3648> A_IWL<3647> A_IWL<3646> A_IWL<3645> A_IWL<3644> A_IWL<3643> A_IWL<3642> A_IWL<3641> A_IWL<3640> A_IWL<3639> A_IWL<3638> A_IWL<3637> A_IWL<3636> A_IWL<3635> A_IWL<3634> A_IWL<3633> A_IWL<3632> A_IWL<3631> A_IWL<3630> A_IWL<3629> A_IWL<3628> A_IWL<3627> A_IWL<3626> A_IWL<3625> A_IWL<3624> A_IWL<3623> A_IWL<3622> A_IWL<3621> A_IWL<3620> A_IWL<3619> A_IWL<3618> A_IWL<3617> A_IWL<3616> A_IWL<3615> A_IWL<3614> A_IWL<3613> A_IWL<3612> A_IWL<3611> A_IWL<3610> A_IWL<3609> A_IWL<3608> A_IWL<3607> A_IWL<3606> A_IWL<3605> A_IWL<3604> A_IWL<3603> A_IWL<3602> A_IWL<3601> A_IWL<3600> A_IWL<3599> A_IWL<3598> A_IWL<3597> A_IWL<3596> A_IWL<3595> A_IWL<3594> A_IWL<3593> A_IWL<3592> A_IWL<3591> A_IWL<3590> A_IWL<3589> A_IWL<3588> A_IWL<3587> A_IWL<3586> A_IWL<3585> A_IWL<3584> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<6> A_BLC<13> A_BLC<12> A_BLC_TOP<13> A_BLC_TOP<12> A_BLT<13> A_BLT<12> A_BLT_TOP<13> A_BLT_TOP<12> A_IWL<3071> A_IWL<3070> A_IWL<3069> A_IWL<3068> A_IWL<3067> A_IWL<3066> A_IWL<3065> A_IWL<3064> A_IWL<3063> A_IWL<3062> A_IWL<3061> A_IWL<3060> A_IWL<3059> A_IWL<3058> A_IWL<3057> A_IWL<3056> A_IWL<3055> A_IWL<3054> A_IWL<3053> A_IWL<3052> A_IWL<3051> A_IWL<3050> A_IWL<3049> A_IWL<3048> A_IWL<3047> A_IWL<3046> A_IWL<3045> A_IWL<3044> A_IWL<3043> A_IWL<3042> A_IWL<3041> A_IWL<3040> A_IWL<3039> A_IWL<3038> A_IWL<3037> A_IWL<3036> A_IWL<3035> A_IWL<3034> A_IWL<3033> A_IWL<3032> A_IWL<3031> A_IWL<3030> A_IWL<3029> A_IWL<3028> A_IWL<3027> A_IWL<3026> A_IWL<3025> A_IWL<3024> A_IWL<3023> A_IWL<3022> A_IWL<3021> A_IWL<3020> A_IWL<3019> A_IWL<3018> A_IWL<3017> A_IWL<3016> A_IWL<3015> A_IWL<3014> A_IWL<3013> A_IWL<3012> A_IWL<3011> A_IWL<3010> A_IWL<3009> A_IWL<3008> A_IWL<3007> A_IWL<3006> A_IWL<3005> A_IWL<3004> A_IWL<3003> A_IWL<3002> A_IWL<3001> A_IWL<3000> A_IWL<2999> A_IWL<2998> A_IWL<2997> A_IWL<2996> A_IWL<2995> A_IWL<2994> A_IWL<2993> A_IWL<2992> A_IWL<2991> A_IWL<2990> A_IWL<2989> A_IWL<2988> A_IWL<2987> A_IWL<2986> A_IWL<2985> A_IWL<2984> A_IWL<2983> A_IWL<2982> A_IWL<2981> A_IWL<2980> A_IWL<2979> A_IWL<2978> A_IWL<2977> A_IWL<2976> A_IWL<2975> A_IWL<2974> A_IWL<2973> A_IWL<2972> A_IWL<2971> A_IWL<2970> A_IWL<2969> A_IWL<2968> A_IWL<2967> A_IWL<2966> A_IWL<2965> A_IWL<2964> A_IWL<2963> A_IWL<2962> A_IWL<2961> A_IWL<2960> A_IWL<2959> A_IWL<2958> A_IWL<2957> A_IWL<2956> A_IWL<2955> A_IWL<2954> A_IWL<2953> A_IWL<2952> A_IWL<2951> A_IWL<2950> A_IWL<2949> A_IWL<2948> A_IWL<2947> A_IWL<2946> A_IWL<2945> A_IWL<2944> A_IWL<2943> A_IWL<2942> A_IWL<2941> A_IWL<2940> A_IWL<2939> A_IWL<2938> A_IWL<2937> A_IWL<2936> A_IWL<2935> A_IWL<2934> A_IWL<2933> A_IWL<2932> A_IWL<2931> A_IWL<2930> A_IWL<2929> A_IWL<2928> A_IWL<2927> A_IWL<2926> A_IWL<2925> A_IWL<2924> A_IWL<2923> A_IWL<2922> A_IWL<2921> A_IWL<2920> A_IWL<2919> A_IWL<2918> A_IWL<2917> A_IWL<2916> A_IWL<2915> A_IWL<2914> A_IWL<2913> A_IWL<2912> A_IWL<2911> A_IWL<2910> A_IWL<2909> A_IWL<2908> A_IWL<2907> A_IWL<2906> A_IWL<2905> A_IWL<2904> A_IWL<2903> A_IWL<2902> A_IWL<2901> A_IWL<2900> A_IWL<2899> A_IWL<2898> A_IWL<2897> A_IWL<2896> A_IWL<2895> A_IWL<2894> A_IWL<2893> A_IWL<2892> A_IWL<2891> A_IWL<2890> A_IWL<2889> A_IWL<2888> A_IWL<2887> A_IWL<2886> A_IWL<2885> A_IWL<2884> A_IWL<2883> A_IWL<2882> A_IWL<2881> A_IWL<2880> A_IWL<2879> A_IWL<2878> A_IWL<2877> A_IWL<2876> A_IWL<2875> A_IWL<2874> A_IWL<2873> A_IWL<2872> A_IWL<2871> A_IWL<2870> A_IWL<2869> A_IWL<2868> A_IWL<2867> A_IWL<2866> A_IWL<2865> A_IWL<2864> A_IWL<2863> A_IWL<2862> A_IWL<2861> A_IWL<2860> A_IWL<2859> A_IWL<2858> A_IWL<2857> A_IWL<2856> A_IWL<2855> A_IWL<2854> A_IWL<2853> A_IWL<2852> A_IWL<2851> A_IWL<2850> A_IWL<2849> A_IWL<2848> A_IWL<2847> A_IWL<2846> A_IWL<2845> A_IWL<2844> A_IWL<2843> A_IWL<2842> A_IWL<2841> A_IWL<2840> A_IWL<2839> A_IWL<2838> A_IWL<2837> A_IWL<2836> A_IWL<2835> A_IWL<2834> A_IWL<2833> A_IWL<2832> A_IWL<2831> A_IWL<2830> A_IWL<2829> A_IWL<2828> A_IWL<2827> A_IWL<2826> A_IWL<2825> A_IWL<2824> A_IWL<2823> A_IWL<2822> A_IWL<2821> A_IWL<2820> A_IWL<2819> A_IWL<2818> A_IWL<2817> A_IWL<2816> A_IWL<2815> A_IWL<2814> A_IWL<2813> A_IWL<2812> A_IWL<2811> A_IWL<2810> A_IWL<2809> A_IWL<2808> A_IWL<2807> A_IWL<2806> A_IWL<2805> A_IWL<2804> A_IWL<2803> A_IWL<2802> A_IWL<2801> A_IWL<2800> A_IWL<2799> A_IWL<2798> A_IWL<2797> A_IWL<2796> A_IWL<2795> A_IWL<2794> A_IWL<2793> A_IWL<2792> A_IWL<2791> A_IWL<2790> A_IWL<2789> A_IWL<2788> A_IWL<2787> A_IWL<2786> A_IWL<2785> A_IWL<2784> A_IWL<2783> A_IWL<2782> A_IWL<2781> A_IWL<2780> A_IWL<2779> A_IWL<2778> A_IWL<2777> A_IWL<2776> A_IWL<2775> A_IWL<2774> A_IWL<2773> A_IWL<2772> A_IWL<2771> A_IWL<2770> A_IWL<2769> A_IWL<2768> A_IWL<2767> A_IWL<2766> A_IWL<2765> A_IWL<2764> A_IWL<2763> A_IWL<2762> A_IWL<2761> A_IWL<2760> A_IWL<2759> A_IWL<2758> A_IWL<2757> A_IWL<2756> A_IWL<2755> A_IWL<2754> A_IWL<2753> A_IWL<2752> A_IWL<2751> A_IWL<2750> A_IWL<2749> A_IWL<2748> A_IWL<2747> A_IWL<2746> A_IWL<2745> A_IWL<2744> A_IWL<2743> A_IWL<2742> A_IWL<2741> A_IWL<2740> A_IWL<2739> A_IWL<2738> A_IWL<2737> A_IWL<2736> A_IWL<2735> A_IWL<2734> A_IWL<2733> A_IWL<2732> A_IWL<2731> A_IWL<2730> A_IWL<2729> A_IWL<2728> A_IWL<2727> A_IWL<2726> A_IWL<2725> A_IWL<2724> A_IWL<2723> A_IWL<2722> A_IWL<2721> A_IWL<2720> A_IWL<2719> A_IWL<2718> A_IWL<2717> A_IWL<2716> A_IWL<2715> A_IWL<2714> A_IWL<2713> A_IWL<2712> A_IWL<2711> A_IWL<2710> A_IWL<2709> A_IWL<2708> A_IWL<2707> A_IWL<2706> A_IWL<2705> A_IWL<2704> A_IWL<2703> A_IWL<2702> A_IWL<2701> A_IWL<2700> A_IWL<2699> A_IWL<2698> A_IWL<2697> A_IWL<2696> A_IWL<2695> A_IWL<2694> A_IWL<2693> A_IWL<2692> A_IWL<2691> A_IWL<2690> A_IWL<2689> A_IWL<2688> A_IWL<2687> A_IWL<2686> A_IWL<2685> A_IWL<2684> A_IWL<2683> A_IWL<2682> A_IWL<2681> A_IWL<2680> A_IWL<2679> A_IWL<2678> A_IWL<2677> A_IWL<2676> A_IWL<2675> A_IWL<2674> A_IWL<2673> A_IWL<2672> A_IWL<2671> A_IWL<2670> A_IWL<2669> A_IWL<2668> A_IWL<2667> A_IWL<2666> A_IWL<2665> A_IWL<2664> A_IWL<2663> A_IWL<2662> A_IWL<2661> A_IWL<2660> A_IWL<2659> A_IWL<2658> A_IWL<2657> A_IWL<2656> A_IWL<2655> A_IWL<2654> A_IWL<2653> A_IWL<2652> A_IWL<2651> A_IWL<2650> A_IWL<2649> A_IWL<2648> A_IWL<2647> A_IWL<2646> A_IWL<2645> A_IWL<2644> A_IWL<2643> A_IWL<2642> A_IWL<2641> A_IWL<2640> A_IWL<2639> A_IWL<2638> A_IWL<2637> A_IWL<2636> A_IWL<2635> A_IWL<2634> A_IWL<2633> A_IWL<2632> A_IWL<2631> A_IWL<2630> A_IWL<2629> A_IWL<2628> A_IWL<2627> A_IWL<2626> A_IWL<2625> A_IWL<2624> A_IWL<2623> A_IWL<2622> A_IWL<2621> A_IWL<2620> A_IWL<2619> A_IWL<2618> A_IWL<2617> A_IWL<2616> A_IWL<2615> A_IWL<2614> A_IWL<2613> A_IWL<2612> A_IWL<2611> A_IWL<2610> A_IWL<2609> A_IWL<2608> A_IWL<2607> A_IWL<2606> A_IWL<2605> A_IWL<2604> A_IWL<2603> A_IWL<2602> A_IWL<2601> A_IWL<2600> A_IWL<2599> A_IWL<2598> A_IWL<2597> A_IWL<2596> A_IWL<2595> A_IWL<2594> A_IWL<2593> A_IWL<2592> A_IWL<2591> A_IWL<2590> A_IWL<2589> A_IWL<2588> A_IWL<2587> A_IWL<2586> A_IWL<2585> A_IWL<2584> A_IWL<2583> A_IWL<2582> A_IWL<2581> A_IWL<2580> A_IWL<2579> A_IWL<2578> A_IWL<2577> A_IWL<2576> A_IWL<2575> A_IWL<2574> A_IWL<2573> A_IWL<2572> A_IWL<2571> A_IWL<2570> A_IWL<2569> A_IWL<2568> A_IWL<2567> A_IWL<2566> A_IWL<2565> A_IWL<2564> A_IWL<2563> A_IWL<2562> A_IWL<2561> A_IWL<2560> A_IWL<3583> A_IWL<3582> A_IWL<3581> A_IWL<3580> A_IWL<3579> A_IWL<3578> A_IWL<3577> A_IWL<3576> A_IWL<3575> A_IWL<3574> A_IWL<3573> A_IWL<3572> A_IWL<3571> A_IWL<3570> A_IWL<3569> A_IWL<3568> A_IWL<3567> A_IWL<3566> A_IWL<3565> A_IWL<3564> A_IWL<3563> A_IWL<3562> A_IWL<3561> A_IWL<3560> A_IWL<3559> A_IWL<3558> A_IWL<3557> A_IWL<3556> A_IWL<3555> A_IWL<3554> A_IWL<3553> A_IWL<3552> A_IWL<3551> A_IWL<3550> A_IWL<3549> A_IWL<3548> A_IWL<3547> A_IWL<3546> A_IWL<3545> A_IWL<3544> A_IWL<3543> A_IWL<3542> A_IWL<3541> A_IWL<3540> A_IWL<3539> A_IWL<3538> A_IWL<3537> A_IWL<3536> A_IWL<3535> A_IWL<3534> A_IWL<3533> A_IWL<3532> A_IWL<3531> A_IWL<3530> A_IWL<3529> A_IWL<3528> A_IWL<3527> A_IWL<3526> A_IWL<3525> A_IWL<3524> A_IWL<3523> A_IWL<3522> A_IWL<3521> A_IWL<3520> A_IWL<3519> A_IWL<3518> A_IWL<3517> A_IWL<3516> A_IWL<3515> A_IWL<3514> A_IWL<3513> A_IWL<3512> A_IWL<3511> A_IWL<3510> A_IWL<3509> A_IWL<3508> A_IWL<3507> A_IWL<3506> A_IWL<3505> A_IWL<3504> A_IWL<3503> A_IWL<3502> A_IWL<3501> A_IWL<3500> A_IWL<3499> A_IWL<3498> A_IWL<3497> A_IWL<3496> A_IWL<3495> A_IWL<3494> A_IWL<3493> A_IWL<3492> A_IWL<3491> A_IWL<3490> A_IWL<3489> A_IWL<3488> A_IWL<3487> A_IWL<3486> A_IWL<3485> A_IWL<3484> A_IWL<3483> A_IWL<3482> A_IWL<3481> A_IWL<3480> A_IWL<3479> A_IWL<3478> A_IWL<3477> A_IWL<3476> A_IWL<3475> A_IWL<3474> A_IWL<3473> A_IWL<3472> A_IWL<3471> A_IWL<3470> A_IWL<3469> A_IWL<3468> A_IWL<3467> A_IWL<3466> A_IWL<3465> A_IWL<3464> A_IWL<3463> A_IWL<3462> A_IWL<3461> A_IWL<3460> A_IWL<3459> A_IWL<3458> A_IWL<3457> A_IWL<3456> A_IWL<3455> A_IWL<3454> A_IWL<3453> A_IWL<3452> A_IWL<3451> A_IWL<3450> A_IWL<3449> A_IWL<3448> A_IWL<3447> A_IWL<3446> A_IWL<3445> A_IWL<3444> A_IWL<3443> A_IWL<3442> A_IWL<3441> A_IWL<3440> A_IWL<3439> A_IWL<3438> A_IWL<3437> A_IWL<3436> A_IWL<3435> A_IWL<3434> A_IWL<3433> A_IWL<3432> A_IWL<3431> A_IWL<3430> A_IWL<3429> A_IWL<3428> A_IWL<3427> A_IWL<3426> A_IWL<3425> A_IWL<3424> A_IWL<3423> A_IWL<3422> A_IWL<3421> A_IWL<3420> A_IWL<3419> A_IWL<3418> A_IWL<3417> A_IWL<3416> A_IWL<3415> A_IWL<3414> A_IWL<3413> A_IWL<3412> A_IWL<3411> A_IWL<3410> A_IWL<3409> A_IWL<3408> A_IWL<3407> A_IWL<3406> A_IWL<3405> A_IWL<3404> A_IWL<3403> A_IWL<3402> A_IWL<3401> A_IWL<3400> A_IWL<3399> A_IWL<3398> A_IWL<3397> A_IWL<3396> A_IWL<3395> A_IWL<3394> A_IWL<3393> A_IWL<3392> A_IWL<3391> A_IWL<3390> A_IWL<3389> A_IWL<3388> A_IWL<3387> A_IWL<3386> A_IWL<3385> A_IWL<3384> A_IWL<3383> A_IWL<3382> A_IWL<3381> A_IWL<3380> A_IWL<3379> A_IWL<3378> A_IWL<3377> A_IWL<3376> A_IWL<3375> A_IWL<3374> A_IWL<3373> A_IWL<3372> A_IWL<3371> A_IWL<3370> A_IWL<3369> A_IWL<3368> A_IWL<3367> A_IWL<3366> A_IWL<3365> A_IWL<3364> A_IWL<3363> A_IWL<3362> A_IWL<3361> A_IWL<3360> A_IWL<3359> A_IWL<3358> A_IWL<3357> A_IWL<3356> A_IWL<3355> A_IWL<3354> A_IWL<3353> A_IWL<3352> A_IWL<3351> A_IWL<3350> A_IWL<3349> A_IWL<3348> A_IWL<3347> A_IWL<3346> A_IWL<3345> A_IWL<3344> A_IWL<3343> A_IWL<3342> A_IWL<3341> A_IWL<3340> A_IWL<3339> A_IWL<3338> A_IWL<3337> A_IWL<3336> A_IWL<3335> A_IWL<3334> A_IWL<3333> A_IWL<3332> A_IWL<3331> A_IWL<3330> A_IWL<3329> A_IWL<3328> A_IWL<3327> A_IWL<3326> A_IWL<3325> A_IWL<3324> A_IWL<3323> A_IWL<3322> A_IWL<3321> A_IWL<3320> A_IWL<3319> A_IWL<3318> A_IWL<3317> A_IWL<3316> A_IWL<3315> A_IWL<3314> A_IWL<3313> A_IWL<3312> A_IWL<3311> A_IWL<3310> A_IWL<3309> A_IWL<3308> A_IWL<3307> A_IWL<3306> A_IWL<3305> A_IWL<3304> A_IWL<3303> A_IWL<3302> A_IWL<3301> A_IWL<3300> A_IWL<3299> A_IWL<3298> A_IWL<3297> A_IWL<3296> A_IWL<3295> A_IWL<3294> A_IWL<3293> A_IWL<3292> A_IWL<3291> A_IWL<3290> A_IWL<3289> A_IWL<3288> A_IWL<3287> A_IWL<3286> A_IWL<3285> A_IWL<3284> A_IWL<3283> A_IWL<3282> A_IWL<3281> A_IWL<3280> A_IWL<3279> A_IWL<3278> A_IWL<3277> A_IWL<3276> A_IWL<3275> A_IWL<3274> A_IWL<3273> A_IWL<3272> A_IWL<3271> A_IWL<3270> A_IWL<3269> A_IWL<3268> A_IWL<3267> A_IWL<3266> A_IWL<3265> A_IWL<3264> A_IWL<3263> A_IWL<3262> A_IWL<3261> A_IWL<3260> A_IWL<3259> A_IWL<3258> A_IWL<3257> A_IWL<3256> A_IWL<3255> A_IWL<3254> A_IWL<3253> A_IWL<3252> A_IWL<3251> A_IWL<3250> A_IWL<3249> A_IWL<3248> A_IWL<3247> A_IWL<3246> A_IWL<3245> A_IWL<3244> A_IWL<3243> A_IWL<3242> A_IWL<3241> A_IWL<3240> A_IWL<3239> A_IWL<3238> A_IWL<3237> A_IWL<3236> A_IWL<3235> A_IWL<3234> A_IWL<3233> A_IWL<3232> A_IWL<3231> A_IWL<3230> A_IWL<3229> A_IWL<3228> A_IWL<3227> A_IWL<3226> A_IWL<3225> A_IWL<3224> A_IWL<3223> A_IWL<3222> A_IWL<3221> A_IWL<3220> A_IWL<3219> A_IWL<3218> A_IWL<3217> A_IWL<3216> A_IWL<3215> A_IWL<3214> A_IWL<3213> A_IWL<3212> A_IWL<3211> A_IWL<3210> A_IWL<3209> A_IWL<3208> A_IWL<3207> A_IWL<3206> A_IWL<3205> A_IWL<3204> A_IWL<3203> A_IWL<3202> A_IWL<3201> A_IWL<3200> A_IWL<3199> A_IWL<3198> A_IWL<3197> A_IWL<3196> A_IWL<3195> A_IWL<3194> A_IWL<3193> A_IWL<3192> A_IWL<3191> A_IWL<3190> A_IWL<3189> A_IWL<3188> A_IWL<3187> A_IWL<3186> A_IWL<3185> A_IWL<3184> A_IWL<3183> A_IWL<3182> A_IWL<3181> A_IWL<3180> A_IWL<3179> A_IWL<3178> A_IWL<3177> A_IWL<3176> A_IWL<3175> A_IWL<3174> A_IWL<3173> A_IWL<3172> A_IWL<3171> A_IWL<3170> A_IWL<3169> A_IWL<3168> A_IWL<3167> A_IWL<3166> A_IWL<3165> A_IWL<3164> A_IWL<3163> A_IWL<3162> A_IWL<3161> A_IWL<3160> A_IWL<3159> A_IWL<3158> A_IWL<3157> A_IWL<3156> A_IWL<3155> A_IWL<3154> A_IWL<3153> A_IWL<3152> A_IWL<3151> A_IWL<3150> A_IWL<3149> A_IWL<3148> A_IWL<3147> A_IWL<3146> A_IWL<3145> A_IWL<3144> A_IWL<3143> A_IWL<3142> A_IWL<3141> A_IWL<3140> A_IWL<3139> A_IWL<3138> A_IWL<3137> A_IWL<3136> A_IWL<3135> A_IWL<3134> A_IWL<3133> A_IWL<3132> A_IWL<3131> A_IWL<3130> A_IWL<3129> A_IWL<3128> A_IWL<3127> A_IWL<3126> A_IWL<3125> A_IWL<3124> A_IWL<3123> A_IWL<3122> A_IWL<3121> A_IWL<3120> A_IWL<3119> A_IWL<3118> A_IWL<3117> A_IWL<3116> A_IWL<3115> A_IWL<3114> A_IWL<3113> A_IWL<3112> A_IWL<3111> A_IWL<3110> A_IWL<3109> A_IWL<3108> A_IWL<3107> A_IWL<3106> A_IWL<3105> A_IWL<3104> A_IWL<3103> A_IWL<3102> A_IWL<3101> A_IWL<3100> A_IWL<3099> A_IWL<3098> A_IWL<3097> A_IWL<3096> A_IWL<3095> A_IWL<3094> A_IWL<3093> A_IWL<3092> A_IWL<3091> A_IWL<3090> A_IWL<3089> A_IWL<3088> A_IWL<3087> A_IWL<3086> A_IWL<3085> A_IWL<3084> A_IWL<3083> A_IWL<3082> A_IWL<3081> A_IWL<3080> A_IWL<3079> A_IWL<3078> A_IWL<3077> A_IWL<3076> A_IWL<3075> A_IWL<3074> A_IWL<3073> A_IWL<3072> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<5> A_BLC<11> A_BLC<10> A_BLC_TOP<11> A_BLC_TOP<10> A_BLT<11> A_BLT<10> A_BLT_TOP<11> A_BLT_TOP<10> A_IWL<2559> A_IWL<2558> A_IWL<2557> A_IWL<2556> A_IWL<2555> A_IWL<2554> A_IWL<2553> A_IWL<2552> A_IWL<2551> A_IWL<2550> A_IWL<2549> A_IWL<2548> A_IWL<2547> A_IWL<2546> A_IWL<2545> A_IWL<2544> A_IWL<2543> A_IWL<2542> A_IWL<2541> A_IWL<2540> A_IWL<2539> A_IWL<2538> A_IWL<2537> A_IWL<2536> A_IWL<2535> A_IWL<2534> A_IWL<2533> A_IWL<2532> A_IWL<2531> A_IWL<2530> A_IWL<2529> A_IWL<2528> A_IWL<2527> A_IWL<2526> A_IWL<2525> A_IWL<2524> A_IWL<2523> A_IWL<2522> A_IWL<2521> A_IWL<2520> A_IWL<2519> A_IWL<2518> A_IWL<2517> A_IWL<2516> A_IWL<2515> A_IWL<2514> A_IWL<2513> A_IWL<2512> A_IWL<2511> A_IWL<2510> A_IWL<2509> A_IWL<2508> A_IWL<2507> A_IWL<2506> A_IWL<2505> A_IWL<2504> A_IWL<2503> A_IWL<2502> A_IWL<2501> A_IWL<2500> A_IWL<2499> A_IWL<2498> A_IWL<2497> A_IWL<2496> A_IWL<2495> A_IWL<2494> A_IWL<2493> A_IWL<2492> A_IWL<2491> A_IWL<2490> A_IWL<2489> A_IWL<2488> A_IWL<2487> A_IWL<2486> A_IWL<2485> A_IWL<2484> A_IWL<2483> A_IWL<2482> A_IWL<2481> A_IWL<2480> A_IWL<2479> A_IWL<2478> A_IWL<2477> A_IWL<2476> A_IWL<2475> A_IWL<2474> A_IWL<2473> A_IWL<2472> A_IWL<2471> A_IWL<2470> A_IWL<2469> A_IWL<2468> A_IWL<2467> A_IWL<2466> A_IWL<2465> A_IWL<2464> A_IWL<2463> A_IWL<2462> A_IWL<2461> A_IWL<2460> A_IWL<2459> A_IWL<2458> A_IWL<2457> A_IWL<2456> A_IWL<2455> A_IWL<2454> A_IWL<2453> A_IWL<2452> A_IWL<2451> A_IWL<2450> A_IWL<2449> A_IWL<2448> A_IWL<2447> A_IWL<2446> A_IWL<2445> A_IWL<2444> A_IWL<2443> A_IWL<2442> A_IWL<2441> A_IWL<2440> A_IWL<2439> A_IWL<2438> A_IWL<2437> A_IWL<2436> A_IWL<2435> A_IWL<2434> A_IWL<2433> A_IWL<2432> A_IWL<2431> A_IWL<2430> A_IWL<2429> A_IWL<2428> A_IWL<2427> A_IWL<2426> A_IWL<2425> A_IWL<2424> A_IWL<2423> A_IWL<2422> A_IWL<2421> A_IWL<2420> A_IWL<2419> A_IWL<2418> A_IWL<2417> A_IWL<2416> A_IWL<2415> A_IWL<2414> A_IWL<2413> A_IWL<2412> A_IWL<2411> A_IWL<2410> A_IWL<2409> A_IWL<2408> A_IWL<2407> A_IWL<2406> A_IWL<2405> A_IWL<2404> A_IWL<2403> A_IWL<2402> A_IWL<2401> A_IWL<2400> A_IWL<2399> A_IWL<2398> A_IWL<2397> A_IWL<2396> A_IWL<2395> A_IWL<2394> A_IWL<2393> A_IWL<2392> A_IWL<2391> A_IWL<2390> A_IWL<2389> A_IWL<2388> A_IWL<2387> A_IWL<2386> A_IWL<2385> A_IWL<2384> A_IWL<2383> A_IWL<2382> A_IWL<2381> A_IWL<2380> A_IWL<2379> A_IWL<2378> A_IWL<2377> A_IWL<2376> A_IWL<2375> A_IWL<2374> A_IWL<2373> A_IWL<2372> A_IWL<2371> A_IWL<2370> A_IWL<2369> A_IWL<2368> A_IWL<2367> A_IWL<2366> A_IWL<2365> A_IWL<2364> A_IWL<2363> A_IWL<2362> A_IWL<2361> A_IWL<2360> A_IWL<2359> A_IWL<2358> A_IWL<2357> A_IWL<2356> A_IWL<2355> A_IWL<2354> A_IWL<2353> A_IWL<2352> A_IWL<2351> A_IWL<2350> A_IWL<2349> A_IWL<2348> A_IWL<2347> A_IWL<2346> A_IWL<2345> A_IWL<2344> A_IWL<2343> A_IWL<2342> A_IWL<2341> A_IWL<2340> A_IWL<2339> A_IWL<2338> A_IWL<2337> A_IWL<2336> A_IWL<2335> A_IWL<2334> A_IWL<2333> A_IWL<2332> A_IWL<2331> A_IWL<2330> A_IWL<2329> A_IWL<2328> A_IWL<2327> A_IWL<2326> A_IWL<2325> A_IWL<2324> A_IWL<2323> A_IWL<2322> A_IWL<2321> A_IWL<2320> A_IWL<2319> A_IWL<2318> A_IWL<2317> A_IWL<2316> A_IWL<2315> A_IWL<2314> A_IWL<2313> A_IWL<2312> A_IWL<2311> A_IWL<2310> A_IWL<2309> A_IWL<2308> A_IWL<2307> A_IWL<2306> A_IWL<2305> A_IWL<2304> A_IWL<2303> A_IWL<2302> A_IWL<2301> A_IWL<2300> A_IWL<2299> A_IWL<2298> A_IWL<2297> A_IWL<2296> A_IWL<2295> A_IWL<2294> A_IWL<2293> A_IWL<2292> A_IWL<2291> A_IWL<2290> A_IWL<2289> A_IWL<2288> A_IWL<2287> A_IWL<2286> A_IWL<2285> A_IWL<2284> A_IWL<2283> A_IWL<2282> A_IWL<2281> A_IWL<2280> A_IWL<2279> A_IWL<2278> A_IWL<2277> A_IWL<2276> A_IWL<2275> A_IWL<2274> A_IWL<2273> A_IWL<2272> A_IWL<2271> A_IWL<2270> A_IWL<2269> A_IWL<2268> A_IWL<2267> A_IWL<2266> A_IWL<2265> A_IWL<2264> A_IWL<2263> A_IWL<2262> A_IWL<2261> A_IWL<2260> A_IWL<2259> A_IWL<2258> A_IWL<2257> A_IWL<2256> A_IWL<2255> A_IWL<2254> A_IWL<2253> A_IWL<2252> A_IWL<2251> A_IWL<2250> A_IWL<2249> A_IWL<2248> A_IWL<2247> A_IWL<2246> A_IWL<2245> A_IWL<2244> A_IWL<2243> A_IWL<2242> A_IWL<2241> A_IWL<2240> A_IWL<2239> A_IWL<2238> A_IWL<2237> A_IWL<2236> A_IWL<2235> A_IWL<2234> A_IWL<2233> A_IWL<2232> A_IWL<2231> A_IWL<2230> A_IWL<2229> A_IWL<2228> A_IWL<2227> A_IWL<2226> A_IWL<2225> A_IWL<2224> A_IWL<2223> A_IWL<2222> A_IWL<2221> A_IWL<2220> A_IWL<2219> A_IWL<2218> A_IWL<2217> A_IWL<2216> A_IWL<2215> A_IWL<2214> A_IWL<2213> A_IWL<2212> A_IWL<2211> A_IWL<2210> A_IWL<2209> A_IWL<2208> A_IWL<2207> A_IWL<2206> A_IWL<2205> A_IWL<2204> A_IWL<2203> A_IWL<2202> A_IWL<2201> A_IWL<2200> A_IWL<2199> A_IWL<2198> A_IWL<2197> A_IWL<2196> A_IWL<2195> A_IWL<2194> A_IWL<2193> A_IWL<2192> A_IWL<2191> A_IWL<2190> A_IWL<2189> A_IWL<2188> A_IWL<2187> A_IWL<2186> A_IWL<2185> A_IWL<2184> A_IWL<2183> A_IWL<2182> A_IWL<2181> A_IWL<2180> A_IWL<2179> A_IWL<2178> A_IWL<2177> A_IWL<2176> A_IWL<2175> A_IWL<2174> A_IWL<2173> A_IWL<2172> A_IWL<2171> A_IWL<2170> A_IWL<2169> A_IWL<2168> A_IWL<2167> A_IWL<2166> A_IWL<2165> A_IWL<2164> A_IWL<2163> A_IWL<2162> A_IWL<2161> A_IWL<2160> A_IWL<2159> A_IWL<2158> A_IWL<2157> A_IWL<2156> A_IWL<2155> A_IWL<2154> A_IWL<2153> A_IWL<2152> A_IWL<2151> A_IWL<2150> A_IWL<2149> A_IWL<2148> A_IWL<2147> A_IWL<2146> A_IWL<2145> A_IWL<2144> A_IWL<2143> A_IWL<2142> A_IWL<2141> A_IWL<2140> A_IWL<2139> A_IWL<2138> A_IWL<2137> A_IWL<2136> A_IWL<2135> A_IWL<2134> A_IWL<2133> A_IWL<2132> A_IWL<2131> A_IWL<2130> A_IWL<2129> A_IWL<2128> A_IWL<2127> A_IWL<2126> A_IWL<2125> A_IWL<2124> A_IWL<2123> A_IWL<2122> A_IWL<2121> A_IWL<2120> A_IWL<2119> A_IWL<2118> A_IWL<2117> A_IWL<2116> A_IWL<2115> A_IWL<2114> A_IWL<2113> A_IWL<2112> A_IWL<2111> A_IWL<2110> A_IWL<2109> A_IWL<2108> A_IWL<2107> A_IWL<2106> A_IWL<2105> A_IWL<2104> A_IWL<2103> A_IWL<2102> A_IWL<2101> A_IWL<2100> A_IWL<2099> A_IWL<2098> A_IWL<2097> A_IWL<2096> A_IWL<2095> A_IWL<2094> A_IWL<2093> A_IWL<2092> A_IWL<2091> A_IWL<2090> A_IWL<2089> A_IWL<2088> A_IWL<2087> A_IWL<2086> A_IWL<2085> A_IWL<2084> A_IWL<2083> A_IWL<2082> A_IWL<2081> A_IWL<2080> A_IWL<2079> A_IWL<2078> A_IWL<2077> A_IWL<2076> A_IWL<2075> A_IWL<2074> A_IWL<2073> A_IWL<2072> A_IWL<2071> A_IWL<2070> A_IWL<2069> A_IWL<2068> A_IWL<2067> A_IWL<2066> A_IWL<2065> A_IWL<2064> A_IWL<2063> A_IWL<2062> A_IWL<2061> A_IWL<2060> A_IWL<2059> A_IWL<2058> A_IWL<2057> A_IWL<2056> A_IWL<2055> A_IWL<2054> A_IWL<2053> A_IWL<2052> A_IWL<2051> A_IWL<2050> A_IWL<2049> A_IWL<2048> A_IWL<3071> A_IWL<3070> A_IWL<3069> A_IWL<3068> A_IWL<3067> A_IWL<3066> A_IWL<3065> A_IWL<3064> A_IWL<3063> A_IWL<3062> A_IWL<3061> A_IWL<3060> A_IWL<3059> A_IWL<3058> A_IWL<3057> A_IWL<3056> A_IWL<3055> A_IWL<3054> A_IWL<3053> A_IWL<3052> A_IWL<3051> A_IWL<3050> A_IWL<3049> A_IWL<3048> A_IWL<3047> A_IWL<3046> A_IWL<3045> A_IWL<3044> A_IWL<3043> A_IWL<3042> A_IWL<3041> A_IWL<3040> A_IWL<3039> A_IWL<3038> A_IWL<3037> A_IWL<3036> A_IWL<3035> A_IWL<3034> A_IWL<3033> A_IWL<3032> A_IWL<3031> A_IWL<3030> A_IWL<3029> A_IWL<3028> A_IWL<3027> A_IWL<3026> A_IWL<3025> A_IWL<3024> A_IWL<3023> A_IWL<3022> A_IWL<3021> A_IWL<3020> A_IWL<3019> A_IWL<3018> A_IWL<3017> A_IWL<3016> A_IWL<3015> A_IWL<3014> A_IWL<3013> A_IWL<3012> A_IWL<3011> A_IWL<3010> A_IWL<3009> A_IWL<3008> A_IWL<3007> A_IWL<3006> A_IWL<3005> A_IWL<3004> A_IWL<3003> A_IWL<3002> A_IWL<3001> A_IWL<3000> A_IWL<2999> A_IWL<2998> A_IWL<2997> A_IWL<2996> A_IWL<2995> A_IWL<2994> A_IWL<2993> A_IWL<2992> A_IWL<2991> A_IWL<2990> A_IWL<2989> A_IWL<2988> A_IWL<2987> A_IWL<2986> A_IWL<2985> A_IWL<2984> A_IWL<2983> A_IWL<2982> A_IWL<2981> A_IWL<2980> A_IWL<2979> A_IWL<2978> A_IWL<2977> A_IWL<2976> A_IWL<2975> A_IWL<2974> A_IWL<2973> A_IWL<2972> A_IWL<2971> A_IWL<2970> A_IWL<2969> A_IWL<2968> A_IWL<2967> A_IWL<2966> A_IWL<2965> A_IWL<2964> A_IWL<2963> A_IWL<2962> A_IWL<2961> A_IWL<2960> A_IWL<2959> A_IWL<2958> A_IWL<2957> A_IWL<2956> A_IWL<2955> A_IWL<2954> A_IWL<2953> A_IWL<2952> A_IWL<2951> A_IWL<2950> A_IWL<2949> A_IWL<2948> A_IWL<2947> A_IWL<2946> A_IWL<2945> A_IWL<2944> A_IWL<2943> A_IWL<2942> A_IWL<2941> A_IWL<2940> A_IWL<2939> A_IWL<2938> A_IWL<2937> A_IWL<2936> A_IWL<2935> A_IWL<2934> A_IWL<2933> A_IWL<2932> A_IWL<2931> A_IWL<2930> A_IWL<2929> A_IWL<2928> A_IWL<2927> A_IWL<2926> A_IWL<2925> A_IWL<2924> A_IWL<2923> A_IWL<2922> A_IWL<2921> A_IWL<2920> A_IWL<2919> A_IWL<2918> A_IWL<2917> A_IWL<2916> A_IWL<2915> A_IWL<2914> A_IWL<2913> A_IWL<2912> A_IWL<2911> A_IWL<2910> A_IWL<2909> A_IWL<2908> A_IWL<2907> A_IWL<2906> A_IWL<2905> A_IWL<2904> A_IWL<2903> A_IWL<2902> A_IWL<2901> A_IWL<2900> A_IWL<2899> A_IWL<2898> A_IWL<2897> A_IWL<2896> A_IWL<2895> A_IWL<2894> A_IWL<2893> A_IWL<2892> A_IWL<2891> A_IWL<2890> A_IWL<2889> A_IWL<2888> A_IWL<2887> A_IWL<2886> A_IWL<2885> A_IWL<2884> A_IWL<2883> A_IWL<2882> A_IWL<2881> A_IWL<2880> A_IWL<2879> A_IWL<2878> A_IWL<2877> A_IWL<2876> A_IWL<2875> A_IWL<2874> A_IWL<2873> A_IWL<2872> A_IWL<2871> A_IWL<2870> A_IWL<2869> A_IWL<2868> A_IWL<2867> A_IWL<2866> A_IWL<2865> A_IWL<2864> A_IWL<2863> A_IWL<2862> A_IWL<2861> A_IWL<2860> A_IWL<2859> A_IWL<2858> A_IWL<2857> A_IWL<2856> A_IWL<2855> A_IWL<2854> A_IWL<2853> A_IWL<2852> A_IWL<2851> A_IWL<2850> A_IWL<2849> A_IWL<2848> A_IWL<2847> A_IWL<2846> A_IWL<2845> A_IWL<2844> A_IWL<2843> A_IWL<2842> A_IWL<2841> A_IWL<2840> A_IWL<2839> A_IWL<2838> A_IWL<2837> A_IWL<2836> A_IWL<2835> A_IWL<2834> A_IWL<2833> A_IWL<2832> A_IWL<2831> A_IWL<2830> A_IWL<2829> A_IWL<2828> A_IWL<2827> A_IWL<2826> A_IWL<2825> A_IWL<2824> A_IWL<2823> A_IWL<2822> A_IWL<2821> A_IWL<2820> A_IWL<2819> A_IWL<2818> A_IWL<2817> A_IWL<2816> A_IWL<2815> A_IWL<2814> A_IWL<2813> A_IWL<2812> A_IWL<2811> A_IWL<2810> A_IWL<2809> A_IWL<2808> A_IWL<2807> A_IWL<2806> A_IWL<2805> A_IWL<2804> A_IWL<2803> A_IWL<2802> A_IWL<2801> A_IWL<2800> A_IWL<2799> A_IWL<2798> A_IWL<2797> A_IWL<2796> A_IWL<2795> A_IWL<2794> A_IWL<2793> A_IWL<2792> A_IWL<2791> A_IWL<2790> A_IWL<2789> A_IWL<2788> A_IWL<2787> A_IWL<2786> A_IWL<2785> A_IWL<2784> A_IWL<2783> A_IWL<2782> A_IWL<2781> A_IWL<2780> A_IWL<2779> A_IWL<2778> A_IWL<2777> A_IWL<2776> A_IWL<2775> A_IWL<2774> A_IWL<2773> A_IWL<2772> A_IWL<2771> A_IWL<2770> A_IWL<2769> A_IWL<2768> A_IWL<2767> A_IWL<2766> A_IWL<2765> A_IWL<2764> A_IWL<2763> A_IWL<2762> A_IWL<2761> A_IWL<2760> A_IWL<2759> A_IWL<2758> A_IWL<2757> A_IWL<2756> A_IWL<2755> A_IWL<2754> A_IWL<2753> A_IWL<2752> A_IWL<2751> A_IWL<2750> A_IWL<2749> A_IWL<2748> A_IWL<2747> A_IWL<2746> A_IWL<2745> A_IWL<2744> A_IWL<2743> A_IWL<2742> A_IWL<2741> A_IWL<2740> A_IWL<2739> A_IWL<2738> A_IWL<2737> A_IWL<2736> A_IWL<2735> A_IWL<2734> A_IWL<2733> A_IWL<2732> A_IWL<2731> A_IWL<2730> A_IWL<2729> A_IWL<2728> A_IWL<2727> A_IWL<2726> A_IWL<2725> A_IWL<2724> A_IWL<2723> A_IWL<2722> A_IWL<2721> A_IWL<2720> A_IWL<2719> A_IWL<2718> A_IWL<2717> A_IWL<2716> A_IWL<2715> A_IWL<2714> A_IWL<2713> A_IWL<2712> A_IWL<2711> A_IWL<2710> A_IWL<2709> A_IWL<2708> A_IWL<2707> A_IWL<2706> A_IWL<2705> A_IWL<2704> A_IWL<2703> A_IWL<2702> A_IWL<2701> A_IWL<2700> A_IWL<2699> A_IWL<2698> A_IWL<2697> A_IWL<2696> A_IWL<2695> A_IWL<2694> A_IWL<2693> A_IWL<2692> A_IWL<2691> A_IWL<2690> A_IWL<2689> A_IWL<2688> A_IWL<2687> A_IWL<2686> A_IWL<2685> A_IWL<2684> A_IWL<2683> A_IWL<2682> A_IWL<2681> A_IWL<2680> A_IWL<2679> A_IWL<2678> A_IWL<2677> A_IWL<2676> A_IWL<2675> A_IWL<2674> A_IWL<2673> A_IWL<2672> A_IWL<2671> A_IWL<2670> A_IWL<2669> A_IWL<2668> A_IWL<2667> A_IWL<2666> A_IWL<2665> A_IWL<2664> A_IWL<2663> A_IWL<2662> A_IWL<2661> A_IWL<2660> A_IWL<2659> A_IWL<2658> A_IWL<2657> A_IWL<2656> A_IWL<2655> A_IWL<2654> A_IWL<2653> A_IWL<2652> A_IWL<2651> A_IWL<2650> A_IWL<2649> A_IWL<2648> A_IWL<2647> A_IWL<2646> A_IWL<2645> A_IWL<2644> A_IWL<2643> A_IWL<2642> A_IWL<2641> A_IWL<2640> A_IWL<2639> A_IWL<2638> A_IWL<2637> A_IWL<2636> A_IWL<2635> A_IWL<2634> A_IWL<2633> A_IWL<2632> A_IWL<2631> A_IWL<2630> A_IWL<2629> A_IWL<2628> A_IWL<2627> A_IWL<2626> A_IWL<2625> A_IWL<2624> A_IWL<2623> A_IWL<2622> A_IWL<2621> A_IWL<2620> A_IWL<2619> A_IWL<2618> A_IWL<2617> A_IWL<2616> A_IWL<2615> A_IWL<2614> A_IWL<2613> A_IWL<2612> A_IWL<2611> A_IWL<2610> A_IWL<2609> A_IWL<2608> A_IWL<2607> A_IWL<2606> A_IWL<2605> A_IWL<2604> A_IWL<2603> A_IWL<2602> A_IWL<2601> A_IWL<2600> A_IWL<2599> A_IWL<2598> A_IWL<2597> A_IWL<2596> A_IWL<2595> A_IWL<2594> A_IWL<2593> A_IWL<2592> A_IWL<2591> A_IWL<2590> A_IWL<2589> A_IWL<2588> A_IWL<2587> A_IWL<2586> A_IWL<2585> A_IWL<2584> A_IWL<2583> A_IWL<2582> A_IWL<2581> A_IWL<2580> A_IWL<2579> A_IWL<2578> A_IWL<2577> A_IWL<2576> A_IWL<2575> A_IWL<2574> A_IWL<2573> A_IWL<2572> A_IWL<2571> A_IWL<2570> A_IWL<2569> A_IWL<2568> A_IWL<2567> A_IWL<2566> A_IWL<2565> A_IWL<2564> A_IWL<2563> A_IWL<2562> A_IWL<2561> A_IWL<2560> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<4> A_BLC<9> A_BLC<8> A_BLC_TOP<9> A_BLC_TOP<8> A_BLT<9> A_BLT<8> A_BLT_TOP<9> A_BLT_TOP<8> A_IWL<2047> A_IWL<2046> A_IWL<2045> A_IWL<2044> A_IWL<2043> A_IWL<2042> A_IWL<2041> A_IWL<2040> A_IWL<2039> A_IWL<2038> A_IWL<2037> A_IWL<2036> A_IWL<2035> A_IWL<2034> A_IWL<2033> A_IWL<2032> A_IWL<2031> A_IWL<2030> A_IWL<2029> A_IWL<2028> A_IWL<2027> A_IWL<2026> A_IWL<2025> A_IWL<2024> A_IWL<2023> A_IWL<2022> A_IWL<2021> A_IWL<2020> A_IWL<2019> A_IWL<2018> A_IWL<2017> A_IWL<2016> A_IWL<2015> A_IWL<2014> A_IWL<2013> A_IWL<2012> A_IWL<2011> A_IWL<2010> A_IWL<2009> A_IWL<2008> A_IWL<2007> A_IWL<2006> A_IWL<2005> A_IWL<2004> A_IWL<2003> A_IWL<2002> A_IWL<2001> A_IWL<2000> A_IWL<1999> A_IWL<1998> A_IWL<1997> A_IWL<1996> A_IWL<1995> A_IWL<1994> A_IWL<1993> A_IWL<1992> A_IWL<1991> A_IWL<1990> A_IWL<1989> A_IWL<1988> A_IWL<1987> A_IWL<1986> A_IWL<1985> A_IWL<1984> A_IWL<1983> A_IWL<1982> A_IWL<1981> A_IWL<1980> A_IWL<1979> A_IWL<1978> A_IWL<1977> A_IWL<1976> A_IWL<1975> A_IWL<1974> A_IWL<1973> A_IWL<1972> A_IWL<1971> A_IWL<1970> A_IWL<1969> A_IWL<1968> A_IWL<1967> A_IWL<1966> A_IWL<1965> A_IWL<1964> A_IWL<1963> A_IWL<1962> A_IWL<1961> A_IWL<1960> A_IWL<1959> A_IWL<1958> A_IWL<1957> A_IWL<1956> A_IWL<1955> A_IWL<1954> A_IWL<1953> A_IWL<1952> A_IWL<1951> A_IWL<1950> A_IWL<1949> A_IWL<1948> A_IWL<1947> A_IWL<1946> A_IWL<1945> A_IWL<1944> A_IWL<1943> A_IWL<1942> A_IWL<1941> A_IWL<1940> A_IWL<1939> A_IWL<1938> A_IWL<1937> A_IWL<1936> A_IWL<1935> A_IWL<1934> A_IWL<1933> A_IWL<1932> A_IWL<1931> A_IWL<1930> A_IWL<1929> A_IWL<1928> A_IWL<1927> A_IWL<1926> A_IWL<1925> A_IWL<1924> A_IWL<1923> A_IWL<1922> A_IWL<1921> A_IWL<1920> A_IWL<1919> A_IWL<1918> A_IWL<1917> A_IWL<1916> A_IWL<1915> A_IWL<1914> A_IWL<1913> A_IWL<1912> A_IWL<1911> A_IWL<1910> A_IWL<1909> A_IWL<1908> A_IWL<1907> A_IWL<1906> A_IWL<1905> A_IWL<1904> A_IWL<1903> A_IWL<1902> A_IWL<1901> A_IWL<1900> A_IWL<1899> A_IWL<1898> A_IWL<1897> A_IWL<1896> A_IWL<1895> A_IWL<1894> A_IWL<1893> A_IWL<1892> A_IWL<1891> A_IWL<1890> A_IWL<1889> A_IWL<1888> A_IWL<1887> A_IWL<1886> A_IWL<1885> A_IWL<1884> A_IWL<1883> A_IWL<1882> A_IWL<1881> A_IWL<1880> A_IWL<1879> A_IWL<1878> A_IWL<1877> A_IWL<1876> A_IWL<1875> A_IWL<1874> A_IWL<1873> A_IWL<1872> A_IWL<1871> A_IWL<1870> A_IWL<1869> A_IWL<1868> A_IWL<1867> A_IWL<1866> A_IWL<1865> A_IWL<1864> A_IWL<1863> A_IWL<1862> A_IWL<1861> A_IWL<1860> A_IWL<1859> A_IWL<1858> A_IWL<1857> A_IWL<1856> A_IWL<1855> A_IWL<1854> A_IWL<1853> A_IWL<1852> A_IWL<1851> A_IWL<1850> A_IWL<1849> A_IWL<1848> A_IWL<1847> A_IWL<1846> A_IWL<1845> A_IWL<1844> A_IWL<1843> A_IWL<1842> A_IWL<1841> A_IWL<1840> A_IWL<1839> A_IWL<1838> A_IWL<1837> A_IWL<1836> A_IWL<1835> A_IWL<1834> A_IWL<1833> A_IWL<1832> A_IWL<1831> A_IWL<1830> A_IWL<1829> A_IWL<1828> A_IWL<1827> A_IWL<1826> A_IWL<1825> A_IWL<1824> A_IWL<1823> A_IWL<1822> A_IWL<1821> A_IWL<1820> A_IWL<1819> A_IWL<1818> A_IWL<1817> A_IWL<1816> A_IWL<1815> A_IWL<1814> A_IWL<1813> A_IWL<1812> A_IWL<1811> A_IWL<1810> A_IWL<1809> A_IWL<1808> A_IWL<1807> A_IWL<1806> A_IWL<1805> A_IWL<1804> A_IWL<1803> A_IWL<1802> A_IWL<1801> A_IWL<1800> A_IWL<1799> A_IWL<1798> A_IWL<1797> A_IWL<1796> A_IWL<1795> A_IWL<1794> A_IWL<1793> A_IWL<1792> A_IWL<1791> A_IWL<1790> A_IWL<1789> A_IWL<1788> A_IWL<1787> A_IWL<1786> A_IWL<1785> A_IWL<1784> A_IWL<1783> A_IWL<1782> A_IWL<1781> A_IWL<1780> A_IWL<1779> A_IWL<1778> A_IWL<1777> A_IWL<1776> A_IWL<1775> A_IWL<1774> A_IWL<1773> A_IWL<1772> A_IWL<1771> A_IWL<1770> A_IWL<1769> A_IWL<1768> A_IWL<1767> A_IWL<1766> A_IWL<1765> A_IWL<1764> A_IWL<1763> A_IWL<1762> A_IWL<1761> A_IWL<1760> A_IWL<1759> A_IWL<1758> A_IWL<1757> A_IWL<1756> A_IWL<1755> A_IWL<1754> A_IWL<1753> A_IWL<1752> A_IWL<1751> A_IWL<1750> A_IWL<1749> A_IWL<1748> A_IWL<1747> A_IWL<1746> A_IWL<1745> A_IWL<1744> A_IWL<1743> A_IWL<1742> A_IWL<1741> A_IWL<1740> A_IWL<1739> A_IWL<1738> A_IWL<1737> A_IWL<1736> A_IWL<1735> A_IWL<1734> A_IWL<1733> A_IWL<1732> A_IWL<1731> A_IWL<1730> A_IWL<1729> A_IWL<1728> A_IWL<1727> A_IWL<1726> A_IWL<1725> A_IWL<1724> A_IWL<1723> A_IWL<1722> A_IWL<1721> A_IWL<1720> A_IWL<1719> A_IWL<1718> A_IWL<1717> A_IWL<1716> A_IWL<1715> A_IWL<1714> A_IWL<1713> A_IWL<1712> A_IWL<1711> A_IWL<1710> A_IWL<1709> A_IWL<1708> A_IWL<1707> A_IWL<1706> A_IWL<1705> A_IWL<1704> A_IWL<1703> A_IWL<1702> A_IWL<1701> A_IWL<1700> A_IWL<1699> A_IWL<1698> A_IWL<1697> A_IWL<1696> A_IWL<1695> A_IWL<1694> A_IWL<1693> A_IWL<1692> A_IWL<1691> A_IWL<1690> A_IWL<1689> A_IWL<1688> A_IWL<1687> A_IWL<1686> A_IWL<1685> A_IWL<1684> A_IWL<1683> A_IWL<1682> A_IWL<1681> A_IWL<1680> A_IWL<1679> A_IWL<1678> A_IWL<1677> A_IWL<1676> A_IWL<1675> A_IWL<1674> A_IWL<1673> A_IWL<1672> A_IWL<1671> A_IWL<1670> A_IWL<1669> A_IWL<1668> A_IWL<1667> A_IWL<1666> A_IWL<1665> A_IWL<1664> A_IWL<1663> A_IWL<1662> A_IWL<1661> A_IWL<1660> A_IWL<1659> A_IWL<1658> A_IWL<1657> A_IWL<1656> A_IWL<1655> A_IWL<1654> A_IWL<1653> A_IWL<1652> A_IWL<1651> A_IWL<1650> A_IWL<1649> A_IWL<1648> A_IWL<1647> A_IWL<1646> A_IWL<1645> A_IWL<1644> A_IWL<1643> A_IWL<1642> A_IWL<1641> A_IWL<1640> A_IWL<1639> A_IWL<1638> A_IWL<1637> A_IWL<1636> A_IWL<1635> A_IWL<1634> A_IWL<1633> A_IWL<1632> A_IWL<1631> A_IWL<1630> A_IWL<1629> A_IWL<1628> A_IWL<1627> A_IWL<1626> A_IWL<1625> A_IWL<1624> A_IWL<1623> A_IWL<1622> A_IWL<1621> A_IWL<1620> A_IWL<1619> A_IWL<1618> A_IWL<1617> A_IWL<1616> A_IWL<1615> A_IWL<1614> A_IWL<1613> A_IWL<1612> A_IWL<1611> A_IWL<1610> A_IWL<1609> A_IWL<1608> A_IWL<1607> A_IWL<1606> A_IWL<1605> A_IWL<1604> A_IWL<1603> A_IWL<1602> A_IWL<1601> A_IWL<1600> A_IWL<1599> A_IWL<1598> A_IWL<1597> A_IWL<1596> A_IWL<1595> A_IWL<1594> A_IWL<1593> A_IWL<1592> A_IWL<1591> A_IWL<1590> A_IWL<1589> A_IWL<1588> A_IWL<1587> A_IWL<1586> A_IWL<1585> A_IWL<1584> A_IWL<1583> A_IWL<1582> A_IWL<1581> A_IWL<1580> A_IWL<1579> A_IWL<1578> A_IWL<1577> A_IWL<1576> A_IWL<1575> A_IWL<1574> A_IWL<1573> A_IWL<1572> A_IWL<1571> A_IWL<1570> A_IWL<1569> A_IWL<1568> A_IWL<1567> A_IWL<1566> A_IWL<1565> A_IWL<1564> A_IWL<1563> A_IWL<1562> A_IWL<1561> A_IWL<1560> A_IWL<1559> A_IWL<1558> A_IWL<1557> A_IWL<1556> A_IWL<1555> A_IWL<1554> A_IWL<1553> A_IWL<1552> A_IWL<1551> A_IWL<1550> A_IWL<1549> A_IWL<1548> A_IWL<1547> A_IWL<1546> A_IWL<1545> A_IWL<1544> A_IWL<1543> A_IWL<1542> A_IWL<1541> A_IWL<1540> A_IWL<1539> A_IWL<1538> A_IWL<1537> A_IWL<1536> A_IWL<2559> A_IWL<2558> A_IWL<2557> A_IWL<2556> A_IWL<2555> A_IWL<2554> A_IWL<2553> A_IWL<2552> A_IWL<2551> A_IWL<2550> A_IWL<2549> A_IWL<2548> A_IWL<2547> A_IWL<2546> A_IWL<2545> A_IWL<2544> A_IWL<2543> A_IWL<2542> A_IWL<2541> A_IWL<2540> A_IWL<2539> A_IWL<2538> A_IWL<2537> A_IWL<2536> A_IWL<2535> A_IWL<2534> A_IWL<2533> A_IWL<2532> A_IWL<2531> A_IWL<2530> A_IWL<2529> A_IWL<2528> A_IWL<2527> A_IWL<2526> A_IWL<2525> A_IWL<2524> A_IWL<2523> A_IWL<2522> A_IWL<2521> A_IWL<2520> A_IWL<2519> A_IWL<2518> A_IWL<2517> A_IWL<2516> A_IWL<2515> A_IWL<2514> A_IWL<2513> A_IWL<2512> A_IWL<2511> A_IWL<2510> A_IWL<2509> A_IWL<2508> A_IWL<2507> A_IWL<2506> A_IWL<2505> A_IWL<2504> A_IWL<2503> A_IWL<2502> A_IWL<2501> A_IWL<2500> A_IWL<2499> A_IWL<2498> A_IWL<2497> A_IWL<2496> A_IWL<2495> A_IWL<2494> A_IWL<2493> A_IWL<2492> A_IWL<2491> A_IWL<2490> A_IWL<2489> A_IWL<2488> A_IWL<2487> A_IWL<2486> A_IWL<2485> A_IWL<2484> A_IWL<2483> A_IWL<2482> A_IWL<2481> A_IWL<2480> A_IWL<2479> A_IWL<2478> A_IWL<2477> A_IWL<2476> A_IWL<2475> A_IWL<2474> A_IWL<2473> A_IWL<2472> A_IWL<2471> A_IWL<2470> A_IWL<2469> A_IWL<2468> A_IWL<2467> A_IWL<2466> A_IWL<2465> A_IWL<2464> A_IWL<2463> A_IWL<2462> A_IWL<2461> A_IWL<2460> A_IWL<2459> A_IWL<2458> A_IWL<2457> A_IWL<2456> A_IWL<2455> A_IWL<2454> A_IWL<2453> A_IWL<2452> A_IWL<2451> A_IWL<2450> A_IWL<2449> A_IWL<2448> A_IWL<2447> A_IWL<2446> A_IWL<2445> A_IWL<2444> A_IWL<2443> A_IWL<2442> A_IWL<2441> A_IWL<2440> A_IWL<2439> A_IWL<2438> A_IWL<2437> A_IWL<2436> A_IWL<2435> A_IWL<2434> A_IWL<2433> A_IWL<2432> A_IWL<2431> A_IWL<2430> A_IWL<2429> A_IWL<2428> A_IWL<2427> A_IWL<2426> A_IWL<2425> A_IWL<2424> A_IWL<2423> A_IWL<2422> A_IWL<2421> A_IWL<2420> A_IWL<2419> A_IWL<2418> A_IWL<2417> A_IWL<2416> A_IWL<2415> A_IWL<2414> A_IWL<2413> A_IWL<2412> A_IWL<2411> A_IWL<2410> A_IWL<2409> A_IWL<2408> A_IWL<2407> A_IWL<2406> A_IWL<2405> A_IWL<2404> A_IWL<2403> A_IWL<2402> A_IWL<2401> A_IWL<2400> A_IWL<2399> A_IWL<2398> A_IWL<2397> A_IWL<2396> A_IWL<2395> A_IWL<2394> A_IWL<2393> A_IWL<2392> A_IWL<2391> A_IWL<2390> A_IWL<2389> A_IWL<2388> A_IWL<2387> A_IWL<2386> A_IWL<2385> A_IWL<2384> A_IWL<2383> A_IWL<2382> A_IWL<2381> A_IWL<2380> A_IWL<2379> A_IWL<2378> A_IWL<2377> A_IWL<2376> A_IWL<2375> A_IWL<2374> A_IWL<2373> A_IWL<2372> A_IWL<2371> A_IWL<2370> A_IWL<2369> A_IWL<2368> A_IWL<2367> A_IWL<2366> A_IWL<2365> A_IWL<2364> A_IWL<2363> A_IWL<2362> A_IWL<2361> A_IWL<2360> A_IWL<2359> A_IWL<2358> A_IWL<2357> A_IWL<2356> A_IWL<2355> A_IWL<2354> A_IWL<2353> A_IWL<2352> A_IWL<2351> A_IWL<2350> A_IWL<2349> A_IWL<2348> A_IWL<2347> A_IWL<2346> A_IWL<2345> A_IWL<2344> A_IWL<2343> A_IWL<2342> A_IWL<2341> A_IWL<2340> A_IWL<2339> A_IWL<2338> A_IWL<2337> A_IWL<2336> A_IWL<2335> A_IWL<2334> A_IWL<2333> A_IWL<2332> A_IWL<2331> A_IWL<2330> A_IWL<2329> A_IWL<2328> A_IWL<2327> A_IWL<2326> A_IWL<2325> A_IWL<2324> A_IWL<2323> A_IWL<2322> A_IWL<2321> A_IWL<2320> A_IWL<2319> A_IWL<2318> A_IWL<2317> A_IWL<2316> A_IWL<2315> A_IWL<2314> A_IWL<2313> A_IWL<2312> A_IWL<2311> A_IWL<2310> A_IWL<2309> A_IWL<2308> A_IWL<2307> A_IWL<2306> A_IWL<2305> A_IWL<2304> A_IWL<2303> A_IWL<2302> A_IWL<2301> A_IWL<2300> A_IWL<2299> A_IWL<2298> A_IWL<2297> A_IWL<2296> A_IWL<2295> A_IWL<2294> A_IWL<2293> A_IWL<2292> A_IWL<2291> A_IWL<2290> A_IWL<2289> A_IWL<2288> A_IWL<2287> A_IWL<2286> A_IWL<2285> A_IWL<2284> A_IWL<2283> A_IWL<2282> A_IWL<2281> A_IWL<2280> A_IWL<2279> A_IWL<2278> A_IWL<2277> A_IWL<2276> A_IWL<2275> A_IWL<2274> A_IWL<2273> A_IWL<2272> A_IWL<2271> A_IWL<2270> A_IWL<2269> A_IWL<2268> A_IWL<2267> A_IWL<2266> A_IWL<2265> A_IWL<2264> A_IWL<2263> A_IWL<2262> A_IWL<2261> A_IWL<2260> A_IWL<2259> A_IWL<2258> A_IWL<2257> A_IWL<2256> A_IWL<2255> A_IWL<2254> A_IWL<2253> A_IWL<2252> A_IWL<2251> A_IWL<2250> A_IWL<2249> A_IWL<2248> A_IWL<2247> A_IWL<2246> A_IWL<2245> A_IWL<2244> A_IWL<2243> A_IWL<2242> A_IWL<2241> A_IWL<2240> A_IWL<2239> A_IWL<2238> A_IWL<2237> A_IWL<2236> A_IWL<2235> A_IWL<2234> A_IWL<2233> A_IWL<2232> A_IWL<2231> A_IWL<2230> A_IWL<2229> A_IWL<2228> A_IWL<2227> A_IWL<2226> A_IWL<2225> A_IWL<2224> A_IWL<2223> A_IWL<2222> A_IWL<2221> A_IWL<2220> A_IWL<2219> A_IWL<2218> A_IWL<2217> A_IWL<2216> A_IWL<2215> A_IWL<2214> A_IWL<2213> A_IWL<2212> A_IWL<2211> A_IWL<2210> A_IWL<2209> A_IWL<2208> A_IWL<2207> A_IWL<2206> A_IWL<2205> A_IWL<2204> A_IWL<2203> A_IWL<2202> A_IWL<2201> A_IWL<2200> A_IWL<2199> A_IWL<2198> A_IWL<2197> A_IWL<2196> A_IWL<2195> A_IWL<2194> A_IWL<2193> A_IWL<2192> A_IWL<2191> A_IWL<2190> A_IWL<2189> A_IWL<2188> A_IWL<2187> A_IWL<2186> A_IWL<2185> A_IWL<2184> A_IWL<2183> A_IWL<2182> A_IWL<2181> A_IWL<2180> A_IWL<2179> A_IWL<2178> A_IWL<2177> A_IWL<2176> A_IWL<2175> A_IWL<2174> A_IWL<2173> A_IWL<2172> A_IWL<2171> A_IWL<2170> A_IWL<2169> A_IWL<2168> A_IWL<2167> A_IWL<2166> A_IWL<2165> A_IWL<2164> A_IWL<2163> A_IWL<2162> A_IWL<2161> A_IWL<2160> A_IWL<2159> A_IWL<2158> A_IWL<2157> A_IWL<2156> A_IWL<2155> A_IWL<2154> A_IWL<2153> A_IWL<2152> A_IWL<2151> A_IWL<2150> A_IWL<2149> A_IWL<2148> A_IWL<2147> A_IWL<2146> A_IWL<2145> A_IWL<2144> A_IWL<2143> A_IWL<2142> A_IWL<2141> A_IWL<2140> A_IWL<2139> A_IWL<2138> A_IWL<2137> A_IWL<2136> A_IWL<2135> A_IWL<2134> A_IWL<2133> A_IWL<2132> A_IWL<2131> A_IWL<2130> A_IWL<2129> A_IWL<2128> A_IWL<2127> A_IWL<2126> A_IWL<2125> A_IWL<2124> A_IWL<2123> A_IWL<2122> A_IWL<2121> A_IWL<2120> A_IWL<2119> A_IWL<2118> A_IWL<2117> A_IWL<2116> A_IWL<2115> A_IWL<2114> A_IWL<2113> A_IWL<2112> A_IWL<2111> A_IWL<2110> A_IWL<2109> A_IWL<2108> A_IWL<2107> A_IWL<2106> A_IWL<2105> A_IWL<2104> A_IWL<2103> A_IWL<2102> A_IWL<2101> A_IWL<2100> A_IWL<2099> A_IWL<2098> A_IWL<2097> A_IWL<2096> A_IWL<2095> A_IWL<2094> A_IWL<2093> A_IWL<2092> A_IWL<2091> A_IWL<2090> A_IWL<2089> A_IWL<2088> A_IWL<2087> A_IWL<2086> A_IWL<2085> A_IWL<2084> A_IWL<2083> A_IWL<2082> A_IWL<2081> A_IWL<2080> A_IWL<2079> A_IWL<2078> A_IWL<2077> A_IWL<2076> A_IWL<2075> A_IWL<2074> A_IWL<2073> A_IWL<2072> A_IWL<2071> A_IWL<2070> A_IWL<2069> A_IWL<2068> A_IWL<2067> A_IWL<2066> A_IWL<2065> A_IWL<2064> A_IWL<2063> A_IWL<2062> A_IWL<2061> A_IWL<2060> A_IWL<2059> A_IWL<2058> A_IWL<2057> A_IWL<2056> A_IWL<2055> A_IWL<2054> A_IWL<2053> A_IWL<2052> A_IWL<2051> A_IWL<2050> A_IWL<2049> A_IWL<2048> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<3> A_BLC<7> A_BLC<6> A_BLC_TOP<7> A_BLC_TOP<6> A_BLT<7> A_BLT<6> A_BLT_TOP<7> A_BLT_TOP<6> A_IWL<1535> A_IWL<1534> A_IWL<1533> A_IWL<1532> A_IWL<1531> A_IWL<1530> A_IWL<1529> A_IWL<1528> A_IWL<1527> A_IWL<1526> A_IWL<1525> A_IWL<1524> A_IWL<1523> A_IWL<1522> A_IWL<1521> A_IWL<1520> A_IWL<1519> A_IWL<1518> A_IWL<1517> A_IWL<1516> A_IWL<1515> A_IWL<1514> A_IWL<1513> A_IWL<1512> A_IWL<1511> A_IWL<1510> A_IWL<1509> A_IWL<1508> A_IWL<1507> A_IWL<1506> A_IWL<1505> A_IWL<1504> A_IWL<1503> A_IWL<1502> A_IWL<1501> A_IWL<1500> A_IWL<1499> A_IWL<1498> A_IWL<1497> A_IWL<1496> A_IWL<1495> A_IWL<1494> A_IWL<1493> A_IWL<1492> A_IWL<1491> A_IWL<1490> A_IWL<1489> A_IWL<1488> A_IWL<1487> A_IWL<1486> A_IWL<1485> A_IWL<1484> A_IWL<1483> A_IWL<1482> A_IWL<1481> A_IWL<1480> A_IWL<1479> A_IWL<1478> A_IWL<1477> A_IWL<1476> A_IWL<1475> A_IWL<1474> A_IWL<1473> A_IWL<1472> A_IWL<1471> A_IWL<1470> A_IWL<1469> A_IWL<1468> A_IWL<1467> A_IWL<1466> A_IWL<1465> A_IWL<1464> A_IWL<1463> A_IWL<1462> A_IWL<1461> A_IWL<1460> A_IWL<1459> A_IWL<1458> A_IWL<1457> A_IWL<1456> A_IWL<1455> A_IWL<1454> A_IWL<1453> A_IWL<1452> A_IWL<1451> A_IWL<1450> A_IWL<1449> A_IWL<1448> A_IWL<1447> A_IWL<1446> A_IWL<1445> A_IWL<1444> A_IWL<1443> A_IWL<1442> A_IWL<1441> A_IWL<1440> A_IWL<1439> A_IWL<1438> A_IWL<1437> A_IWL<1436> A_IWL<1435> A_IWL<1434> A_IWL<1433> A_IWL<1432> A_IWL<1431> A_IWL<1430> A_IWL<1429> A_IWL<1428> A_IWL<1427> A_IWL<1426> A_IWL<1425> A_IWL<1424> A_IWL<1423> A_IWL<1422> A_IWL<1421> A_IWL<1420> A_IWL<1419> A_IWL<1418> A_IWL<1417> A_IWL<1416> A_IWL<1415> A_IWL<1414> A_IWL<1413> A_IWL<1412> A_IWL<1411> A_IWL<1410> A_IWL<1409> A_IWL<1408> A_IWL<1407> A_IWL<1406> A_IWL<1405> A_IWL<1404> A_IWL<1403> A_IWL<1402> A_IWL<1401> A_IWL<1400> A_IWL<1399> A_IWL<1398> A_IWL<1397> A_IWL<1396> A_IWL<1395> A_IWL<1394> A_IWL<1393> A_IWL<1392> A_IWL<1391> A_IWL<1390> A_IWL<1389> A_IWL<1388> A_IWL<1387> A_IWL<1386> A_IWL<1385> A_IWL<1384> A_IWL<1383> A_IWL<1382> A_IWL<1381> A_IWL<1380> A_IWL<1379> A_IWL<1378> A_IWL<1377> A_IWL<1376> A_IWL<1375> A_IWL<1374> A_IWL<1373> A_IWL<1372> A_IWL<1371> A_IWL<1370> A_IWL<1369> A_IWL<1368> A_IWL<1367> A_IWL<1366> A_IWL<1365> A_IWL<1364> A_IWL<1363> A_IWL<1362> A_IWL<1361> A_IWL<1360> A_IWL<1359> A_IWL<1358> A_IWL<1357> A_IWL<1356> A_IWL<1355> A_IWL<1354> A_IWL<1353> A_IWL<1352> A_IWL<1351> A_IWL<1350> A_IWL<1349> A_IWL<1348> A_IWL<1347> A_IWL<1346> A_IWL<1345> A_IWL<1344> A_IWL<1343> A_IWL<1342> A_IWL<1341> A_IWL<1340> A_IWL<1339> A_IWL<1338> A_IWL<1337> A_IWL<1336> A_IWL<1335> A_IWL<1334> A_IWL<1333> A_IWL<1332> A_IWL<1331> A_IWL<1330> A_IWL<1329> A_IWL<1328> A_IWL<1327> A_IWL<1326> A_IWL<1325> A_IWL<1324> A_IWL<1323> A_IWL<1322> A_IWL<1321> A_IWL<1320> A_IWL<1319> A_IWL<1318> A_IWL<1317> A_IWL<1316> A_IWL<1315> A_IWL<1314> A_IWL<1313> A_IWL<1312> A_IWL<1311> A_IWL<1310> A_IWL<1309> A_IWL<1308> A_IWL<1307> A_IWL<1306> A_IWL<1305> A_IWL<1304> A_IWL<1303> A_IWL<1302> A_IWL<1301> A_IWL<1300> A_IWL<1299> A_IWL<1298> A_IWL<1297> A_IWL<1296> A_IWL<1295> A_IWL<1294> A_IWL<1293> A_IWL<1292> A_IWL<1291> A_IWL<1290> A_IWL<1289> A_IWL<1288> A_IWL<1287> A_IWL<1286> A_IWL<1285> A_IWL<1284> A_IWL<1283> A_IWL<1282> A_IWL<1281> A_IWL<1280> A_IWL<1279> A_IWL<1278> A_IWL<1277> A_IWL<1276> A_IWL<1275> A_IWL<1274> A_IWL<1273> A_IWL<1272> A_IWL<1271> A_IWL<1270> A_IWL<1269> A_IWL<1268> A_IWL<1267> A_IWL<1266> A_IWL<1265> A_IWL<1264> A_IWL<1263> A_IWL<1262> A_IWL<1261> A_IWL<1260> A_IWL<1259> A_IWL<1258> A_IWL<1257> A_IWL<1256> A_IWL<1255> A_IWL<1254> A_IWL<1253> A_IWL<1252> A_IWL<1251> A_IWL<1250> A_IWL<1249> A_IWL<1248> A_IWL<1247> A_IWL<1246> A_IWL<1245> A_IWL<1244> A_IWL<1243> A_IWL<1242> A_IWL<1241> A_IWL<1240> A_IWL<1239> A_IWL<1238> A_IWL<1237> A_IWL<1236> A_IWL<1235> A_IWL<1234> A_IWL<1233> A_IWL<1232> A_IWL<1231> A_IWL<1230> A_IWL<1229> A_IWL<1228> A_IWL<1227> A_IWL<1226> A_IWL<1225> A_IWL<1224> A_IWL<1223> A_IWL<1222> A_IWL<1221> A_IWL<1220> A_IWL<1219> A_IWL<1218> A_IWL<1217> A_IWL<1216> A_IWL<1215> A_IWL<1214> A_IWL<1213> A_IWL<1212> A_IWL<1211> A_IWL<1210> A_IWL<1209> A_IWL<1208> A_IWL<1207> A_IWL<1206> A_IWL<1205> A_IWL<1204> A_IWL<1203> A_IWL<1202> A_IWL<1201> A_IWL<1200> A_IWL<1199> A_IWL<1198> A_IWL<1197> A_IWL<1196> A_IWL<1195> A_IWL<1194> A_IWL<1193> A_IWL<1192> A_IWL<1191> A_IWL<1190> A_IWL<1189> A_IWL<1188> A_IWL<1187> A_IWL<1186> A_IWL<1185> A_IWL<1184> A_IWL<1183> A_IWL<1182> A_IWL<1181> A_IWL<1180> A_IWL<1179> A_IWL<1178> A_IWL<1177> A_IWL<1176> A_IWL<1175> A_IWL<1174> A_IWL<1173> A_IWL<1172> A_IWL<1171> A_IWL<1170> A_IWL<1169> A_IWL<1168> A_IWL<1167> A_IWL<1166> A_IWL<1165> A_IWL<1164> A_IWL<1163> A_IWL<1162> A_IWL<1161> A_IWL<1160> A_IWL<1159> A_IWL<1158> A_IWL<1157> A_IWL<1156> A_IWL<1155> A_IWL<1154> A_IWL<1153> A_IWL<1152> A_IWL<1151> A_IWL<1150> A_IWL<1149> A_IWL<1148> A_IWL<1147> A_IWL<1146> A_IWL<1145> A_IWL<1144> A_IWL<1143> A_IWL<1142> A_IWL<1141> A_IWL<1140> A_IWL<1139> A_IWL<1138> A_IWL<1137> A_IWL<1136> A_IWL<1135> A_IWL<1134> A_IWL<1133> A_IWL<1132> A_IWL<1131> A_IWL<1130> A_IWL<1129> A_IWL<1128> A_IWL<1127> A_IWL<1126> A_IWL<1125> A_IWL<1124> A_IWL<1123> A_IWL<1122> A_IWL<1121> A_IWL<1120> A_IWL<1119> A_IWL<1118> A_IWL<1117> A_IWL<1116> A_IWL<1115> A_IWL<1114> A_IWL<1113> A_IWL<1112> A_IWL<1111> A_IWL<1110> A_IWL<1109> A_IWL<1108> A_IWL<1107> A_IWL<1106> A_IWL<1105> A_IWL<1104> A_IWL<1103> A_IWL<1102> A_IWL<1101> A_IWL<1100> A_IWL<1099> A_IWL<1098> A_IWL<1097> A_IWL<1096> A_IWL<1095> A_IWL<1094> A_IWL<1093> A_IWL<1092> A_IWL<1091> A_IWL<1090> A_IWL<1089> A_IWL<1088> A_IWL<1087> A_IWL<1086> A_IWL<1085> A_IWL<1084> A_IWL<1083> A_IWL<1082> A_IWL<1081> A_IWL<1080> A_IWL<1079> A_IWL<1078> A_IWL<1077> A_IWL<1076> A_IWL<1075> A_IWL<1074> A_IWL<1073> A_IWL<1072> A_IWL<1071> A_IWL<1070> A_IWL<1069> A_IWL<1068> A_IWL<1067> A_IWL<1066> A_IWL<1065> A_IWL<1064> A_IWL<1063> A_IWL<1062> A_IWL<1061> A_IWL<1060> A_IWL<1059> A_IWL<1058> A_IWL<1057> A_IWL<1056> A_IWL<1055> A_IWL<1054> A_IWL<1053> A_IWL<1052> A_IWL<1051> A_IWL<1050> A_IWL<1049> A_IWL<1048> A_IWL<1047> A_IWL<1046> A_IWL<1045> A_IWL<1044> A_IWL<1043> A_IWL<1042> A_IWL<1041> A_IWL<1040> A_IWL<1039> A_IWL<1038> A_IWL<1037> A_IWL<1036> A_IWL<1035> A_IWL<1034> A_IWL<1033> A_IWL<1032> A_IWL<1031> A_IWL<1030> A_IWL<1029> A_IWL<1028> A_IWL<1027> A_IWL<1026> A_IWL<1025> A_IWL<1024> A_IWL<2047> A_IWL<2046> A_IWL<2045> A_IWL<2044> A_IWL<2043> A_IWL<2042> A_IWL<2041> A_IWL<2040> A_IWL<2039> A_IWL<2038> A_IWL<2037> A_IWL<2036> A_IWL<2035> A_IWL<2034> A_IWL<2033> A_IWL<2032> A_IWL<2031> A_IWL<2030> A_IWL<2029> A_IWL<2028> A_IWL<2027> A_IWL<2026> A_IWL<2025> A_IWL<2024> A_IWL<2023> A_IWL<2022> A_IWL<2021> A_IWL<2020> A_IWL<2019> A_IWL<2018> A_IWL<2017> A_IWL<2016> A_IWL<2015> A_IWL<2014> A_IWL<2013> A_IWL<2012> A_IWL<2011> A_IWL<2010> A_IWL<2009> A_IWL<2008> A_IWL<2007> A_IWL<2006> A_IWL<2005> A_IWL<2004> A_IWL<2003> A_IWL<2002> A_IWL<2001> A_IWL<2000> A_IWL<1999> A_IWL<1998> A_IWL<1997> A_IWL<1996> A_IWL<1995> A_IWL<1994> A_IWL<1993> A_IWL<1992> A_IWL<1991> A_IWL<1990> A_IWL<1989> A_IWL<1988> A_IWL<1987> A_IWL<1986> A_IWL<1985> A_IWL<1984> A_IWL<1983> A_IWL<1982> A_IWL<1981> A_IWL<1980> A_IWL<1979> A_IWL<1978> A_IWL<1977> A_IWL<1976> A_IWL<1975> A_IWL<1974> A_IWL<1973> A_IWL<1972> A_IWL<1971> A_IWL<1970> A_IWL<1969> A_IWL<1968> A_IWL<1967> A_IWL<1966> A_IWL<1965> A_IWL<1964> A_IWL<1963> A_IWL<1962> A_IWL<1961> A_IWL<1960> A_IWL<1959> A_IWL<1958> A_IWL<1957> A_IWL<1956> A_IWL<1955> A_IWL<1954> A_IWL<1953> A_IWL<1952> A_IWL<1951> A_IWL<1950> A_IWL<1949> A_IWL<1948> A_IWL<1947> A_IWL<1946> A_IWL<1945> A_IWL<1944> A_IWL<1943> A_IWL<1942> A_IWL<1941> A_IWL<1940> A_IWL<1939> A_IWL<1938> A_IWL<1937> A_IWL<1936> A_IWL<1935> A_IWL<1934> A_IWL<1933> A_IWL<1932> A_IWL<1931> A_IWL<1930> A_IWL<1929> A_IWL<1928> A_IWL<1927> A_IWL<1926> A_IWL<1925> A_IWL<1924> A_IWL<1923> A_IWL<1922> A_IWL<1921> A_IWL<1920> A_IWL<1919> A_IWL<1918> A_IWL<1917> A_IWL<1916> A_IWL<1915> A_IWL<1914> A_IWL<1913> A_IWL<1912> A_IWL<1911> A_IWL<1910> A_IWL<1909> A_IWL<1908> A_IWL<1907> A_IWL<1906> A_IWL<1905> A_IWL<1904> A_IWL<1903> A_IWL<1902> A_IWL<1901> A_IWL<1900> A_IWL<1899> A_IWL<1898> A_IWL<1897> A_IWL<1896> A_IWL<1895> A_IWL<1894> A_IWL<1893> A_IWL<1892> A_IWL<1891> A_IWL<1890> A_IWL<1889> A_IWL<1888> A_IWL<1887> A_IWL<1886> A_IWL<1885> A_IWL<1884> A_IWL<1883> A_IWL<1882> A_IWL<1881> A_IWL<1880> A_IWL<1879> A_IWL<1878> A_IWL<1877> A_IWL<1876> A_IWL<1875> A_IWL<1874> A_IWL<1873> A_IWL<1872> A_IWL<1871> A_IWL<1870> A_IWL<1869> A_IWL<1868> A_IWL<1867> A_IWL<1866> A_IWL<1865> A_IWL<1864> A_IWL<1863> A_IWL<1862> A_IWL<1861> A_IWL<1860> A_IWL<1859> A_IWL<1858> A_IWL<1857> A_IWL<1856> A_IWL<1855> A_IWL<1854> A_IWL<1853> A_IWL<1852> A_IWL<1851> A_IWL<1850> A_IWL<1849> A_IWL<1848> A_IWL<1847> A_IWL<1846> A_IWL<1845> A_IWL<1844> A_IWL<1843> A_IWL<1842> A_IWL<1841> A_IWL<1840> A_IWL<1839> A_IWL<1838> A_IWL<1837> A_IWL<1836> A_IWL<1835> A_IWL<1834> A_IWL<1833> A_IWL<1832> A_IWL<1831> A_IWL<1830> A_IWL<1829> A_IWL<1828> A_IWL<1827> A_IWL<1826> A_IWL<1825> A_IWL<1824> A_IWL<1823> A_IWL<1822> A_IWL<1821> A_IWL<1820> A_IWL<1819> A_IWL<1818> A_IWL<1817> A_IWL<1816> A_IWL<1815> A_IWL<1814> A_IWL<1813> A_IWL<1812> A_IWL<1811> A_IWL<1810> A_IWL<1809> A_IWL<1808> A_IWL<1807> A_IWL<1806> A_IWL<1805> A_IWL<1804> A_IWL<1803> A_IWL<1802> A_IWL<1801> A_IWL<1800> A_IWL<1799> A_IWL<1798> A_IWL<1797> A_IWL<1796> A_IWL<1795> A_IWL<1794> A_IWL<1793> A_IWL<1792> A_IWL<1791> A_IWL<1790> A_IWL<1789> A_IWL<1788> A_IWL<1787> A_IWL<1786> A_IWL<1785> A_IWL<1784> A_IWL<1783> A_IWL<1782> A_IWL<1781> A_IWL<1780> A_IWL<1779> A_IWL<1778> A_IWL<1777> A_IWL<1776> A_IWL<1775> A_IWL<1774> A_IWL<1773> A_IWL<1772> A_IWL<1771> A_IWL<1770> A_IWL<1769> A_IWL<1768> A_IWL<1767> A_IWL<1766> A_IWL<1765> A_IWL<1764> A_IWL<1763> A_IWL<1762> A_IWL<1761> A_IWL<1760> A_IWL<1759> A_IWL<1758> A_IWL<1757> A_IWL<1756> A_IWL<1755> A_IWL<1754> A_IWL<1753> A_IWL<1752> A_IWL<1751> A_IWL<1750> A_IWL<1749> A_IWL<1748> A_IWL<1747> A_IWL<1746> A_IWL<1745> A_IWL<1744> A_IWL<1743> A_IWL<1742> A_IWL<1741> A_IWL<1740> A_IWL<1739> A_IWL<1738> A_IWL<1737> A_IWL<1736> A_IWL<1735> A_IWL<1734> A_IWL<1733> A_IWL<1732> A_IWL<1731> A_IWL<1730> A_IWL<1729> A_IWL<1728> A_IWL<1727> A_IWL<1726> A_IWL<1725> A_IWL<1724> A_IWL<1723> A_IWL<1722> A_IWL<1721> A_IWL<1720> A_IWL<1719> A_IWL<1718> A_IWL<1717> A_IWL<1716> A_IWL<1715> A_IWL<1714> A_IWL<1713> A_IWL<1712> A_IWL<1711> A_IWL<1710> A_IWL<1709> A_IWL<1708> A_IWL<1707> A_IWL<1706> A_IWL<1705> A_IWL<1704> A_IWL<1703> A_IWL<1702> A_IWL<1701> A_IWL<1700> A_IWL<1699> A_IWL<1698> A_IWL<1697> A_IWL<1696> A_IWL<1695> A_IWL<1694> A_IWL<1693> A_IWL<1692> A_IWL<1691> A_IWL<1690> A_IWL<1689> A_IWL<1688> A_IWL<1687> A_IWL<1686> A_IWL<1685> A_IWL<1684> A_IWL<1683> A_IWL<1682> A_IWL<1681> A_IWL<1680> A_IWL<1679> A_IWL<1678> A_IWL<1677> A_IWL<1676> A_IWL<1675> A_IWL<1674> A_IWL<1673> A_IWL<1672> A_IWL<1671> A_IWL<1670> A_IWL<1669> A_IWL<1668> A_IWL<1667> A_IWL<1666> A_IWL<1665> A_IWL<1664> A_IWL<1663> A_IWL<1662> A_IWL<1661> A_IWL<1660> A_IWL<1659> A_IWL<1658> A_IWL<1657> A_IWL<1656> A_IWL<1655> A_IWL<1654> A_IWL<1653> A_IWL<1652> A_IWL<1651> A_IWL<1650> A_IWL<1649> A_IWL<1648> A_IWL<1647> A_IWL<1646> A_IWL<1645> A_IWL<1644> A_IWL<1643> A_IWL<1642> A_IWL<1641> A_IWL<1640> A_IWL<1639> A_IWL<1638> A_IWL<1637> A_IWL<1636> A_IWL<1635> A_IWL<1634> A_IWL<1633> A_IWL<1632> A_IWL<1631> A_IWL<1630> A_IWL<1629> A_IWL<1628> A_IWL<1627> A_IWL<1626> A_IWL<1625> A_IWL<1624> A_IWL<1623> A_IWL<1622> A_IWL<1621> A_IWL<1620> A_IWL<1619> A_IWL<1618> A_IWL<1617> A_IWL<1616> A_IWL<1615> A_IWL<1614> A_IWL<1613> A_IWL<1612> A_IWL<1611> A_IWL<1610> A_IWL<1609> A_IWL<1608> A_IWL<1607> A_IWL<1606> A_IWL<1605> A_IWL<1604> A_IWL<1603> A_IWL<1602> A_IWL<1601> A_IWL<1600> A_IWL<1599> A_IWL<1598> A_IWL<1597> A_IWL<1596> A_IWL<1595> A_IWL<1594> A_IWL<1593> A_IWL<1592> A_IWL<1591> A_IWL<1590> A_IWL<1589> A_IWL<1588> A_IWL<1587> A_IWL<1586> A_IWL<1585> A_IWL<1584> A_IWL<1583> A_IWL<1582> A_IWL<1581> A_IWL<1580> A_IWL<1579> A_IWL<1578> A_IWL<1577> A_IWL<1576> A_IWL<1575> A_IWL<1574> A_IWL<1573> A_IWL<1572> A_IWL<1571> A_IWL<1570> A_IWL<1569> A_IWL<1568> A_IWL<1567> A_IWL<1566> A_IWL<1565> A_IWL<1564> A_IWL<1563> A_IWL<1562> A_IWL<1561> A_IWL<1560> A_IWL<1559> A_IWL<1558> A_IWL<1557> A_IWL<1556> A_IWL<1555> A_IWL<1554> A_IWL<1553> A_IWL<1552> A_IWL<1551> A_IWL<1550> A_IWL<1549> A_IWL<1548> A_IWL<1547> A_IWL<1546> A_IWL<1545> A_IWL<1544> A_IWL<1543> A_IWL<1542> A_IWL<1541> A_IWL<1540> A_IWL<1539> A_IWL<1538> A_IWL<1537> A_IWL<1536> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<2> A_BLC<5> A_BLC<4> A_BLC_TOP<5> A_BLC_TOP<4> A_BLT<5> A_BLT<4> A_BLT_TOP<5> A_BLT_TOP<4> A_IWL<1023> A_IWL<1022> A_IWL<1021> A_IWL<1020> A_IWL<1019> A_IWL<1018> A_IWL<1017> A_IWL<1016> A_IWL<1015> A_IWL<1014> A_IWL<1013> A_IWL<1012> A_IWL<1011> A_IWL<1010> A_IWL<1009> A_IWL<1008> A_IWL<1007> A_IWL<1006> A_IWL<1005> A_IWL<1004> A_IWL<1003> A_IWL<1002> A_IWL<1001> A_IWL<1000> A_IWL<999> A_IWL<998> A_IWL<997> A_IWL<996> A_IWL<995> A_IWL<994> A_IWL<993> A_IWL<992> A_IWL<991> A_IWL<990> A_IWL<989> A_IWL<988> A_IWL<987> A_IWL<986> A_IWL<985> A_IWL<984> A_IWL<983> A_IWL<982> A_IWL<981> A_IWL<980> A_IWL<979> A_IWL<978> A_IWL<977> A_IWL<976> A_IWL<975> A_IWL<974> A_IWL<973> A_IWL<972> A_IWL<971> A_IWL<970> A_IWL<969> A_IWL<968> A_IWL<967> A_IWL<966> A_IWL<965> A_IWL<964> A_IWL<963> A_IWL<962> A_IWL<961> A_IWL<960> A_IWL<959> A_IWL<958> A_IWL<957> A_IWL<956> A_IWL<955> A_IWL<954> A_IWL<953> A_IWL<952> A_IWL<951> A_IWL<950> A_IWL<949> A_IWL<948> A_IWL<947> A_IWL<946> A_IWL<945> A_IWL<944> A_IWL<943> A_IWL<942> A_IWL<941> A_IWL<940> A_IWL<939> A_IWL<938> A_IWL<937> A_IWL<936> A_IWL<935> A_IWL<934> A_IWL<933> A_IWL<932> A_IWL<931> A_IWL<930> A_IWL<929> A_IWL<928> A_IWL<927> A_IWL<926> A_IWL<925> A_IWL<924> A_IWL<923> A_IWL<922> A_IWL<921> A_IWL<920> A_IWL<919> A_IWL<918> A_IWL<917> A_IWL<916> A_IWL<915> A_IWL<914> A_IWL<913> A_IWL<912> A_IWL<911> A_IWL<910> A_IWL<909> A_IWL<908> A_IWL<907> A_IWL<906> A_IWL<905> A_IWL<904> A_IWL<903> A_IWL<902> A_IWL<901> A_IWL<900> A_IWL<899> A_IWL<898> A_IWL<897> A_IWL<896> A_IWL<895> A_IWL<894> A_IWL<893> A_IWL<892> A_IWL<891> A_IWL<890> A_IWL<889> A_IWL<888> A_IWL<887> A_IWL<886> A_IWL<885> A_IWL<884> A_IWL<883> A_IWL<882> A_IWL<881> A_IWL<880> A_IWL<879> A_IWL<878> A_IWL<877> A_IWL<876> A_IWL<875> A_IWL<874> A_IWL<873> A_IWL<872> A_IWL<871> A_IWL<870> A_IWL<869> A_IWL<868> A_IWL<867> A_IWL<866> A_IWL<865> A_IWL<864> A_IWL<863> A_IWL<862> A_IWL<861> A_IWL<860> A_IWL<859> A_IWL<858> A_IWL<857> A_IWL<856> A_IWL<855> A_IWL<854> A_IWL<853> A_IWL<852> A_IWL<851> A_IWL<850> A_IWL<849> A_IWL<848> A_IWL<847> A_IWL<846> A_IWL<845> A_IWL<844> A_IWL<843> A_IWL<842> A_IWL<841> A_IWL<840> A_IWL<839> A_IWL<838> A_IWL<837> A_IWL<836> A_IWL<835> A_IWL<834> A_IWL<833> A_IWL<832> A_IWL<831> A_IWL<830> A_IWL<829> A_IWL<828> A_IWL<827> A_IWL<826> A_IWL<825> A_IWL<824> A_IWL<823> A_IWL<822> A_IWL<821> A_IWL<820> A_IWL<819> A_IWL<818> A_IWL<817> A_IWL<816> A_IWL<815> A_IWL<814> A_IWL<813> A_IWL<812> A_IWL<811> A_IWL<810> A_IWL<809> A_IWL<808> A_IWL<807> A_IWL<806> A_IWL<805> A_IWL<804> A_IWL<803> A_IWL<802> A_IWL<801> A_IWL<800> A_IWL<799> A_IWL<798> A_IWL<797> A_IWL<796> A_IWL<795> A_IWL<794> A_IWL<793> A_IWL<792> A_IWL<791> A_IWL<790> A_IWL<789> A_IWL<788> A_IWL<787> A_IWL<786> A_IWL<785> A_IWL<784> A_IWL<783> A_IWL<782> A_IWL<781> A_IWL<780> A_IWL<779> A_IWL<778> A_IWL<777> A_IWL<776> A_IWL<775> A_IWL<774> A_IWL<773> A_IWL<772> A_IWL<771> A_IWL<770> A_IWL<769> A_IWL<768> A_IWL<767> A_IWL<766> A_IWL<765> A_IWL<764> A_IWL<763> A_IWL<762> A_IWL<761> A_IWL<760> A_IWL<759> A_IWL<758> A_IWL<757> A_IWL<756> A_IWL<755> A_IWL<754> A_IWL<753> A_IWL<752> A_IWL<751> A_IWL<750> A_IWL<749> A_IWL<748> A_IWL<747> A_IWL<746> A_IWL<745> A_IWL<744> A_IWL<743> A_IWL<742> A_IWL<741> A_IWL<740> A_IWL<739> A_IWL<738> A_IWL<737> A_IWL<736> A_IWL<735> A_IWL<734> A_IWL<733> A_IWL<732> A_IWL<731> A_IWL<730> A_IWL<729> A_IWL<728> A_IWL<727> A_IWL<726> A_IWL<725> A_IWL<724> A_IWL<723> A_IWL<722> A_IWL<721> A_IWL<720> A_IWL<719> A_IWL<718> A_IWL<717> A_IWL<716> A_IWL<715> A_IWL<714> A_IWL<713> A_IWL<712> A_IWL<711> A_IWL<710> A_IWL<709> A_IWL<708> A_IWL<707> A_IWL<706> A_IWL<705> A_IWL<704> A_IWL<703> A_IWL<702> A_IWL<701> A_IWL<700> A_IWL<699> A_IWL<698> A_IWL<697> A_IWL<696> A_IWL<695> A_IWL<694> A_IWL<693> A_IWL<692> A_IWL<691> A_IWL<690> A_IWL<689> A_IWL<688> A_IWL<687> A_IWL<686> A_IWL<685> A_IWL<684> A_IWL<683> A_IWL<682> A_IWL<681> A_IWL<680> A_IWL<679> A_IWL<678> A_IWL<677> A_IWL<676> A_IWL<675> A_IWL<674> A_IWL<673> A_IWL<672> A_IWL<671> A_IWL<670> A_IWL<669> A_IWL<668> A_IWL<667> A_IWL<666> A_IWL<665> A_IWL<664> A_IWL<663> A_IWL<662> A_IWL<661> A_IWL<660> A_IWL<659> A_IWL<658> A_IWL<657> A_IWL<656> A_IWL<655> A_IWL<654> A_IWL<653> A_IWL<652> A_IWL<651> A_IWL<650> A_IWL<649> A_IWL<648> A_IWL<647> A_IWL<646> A_IWL<645> A_IWL<644> A_IWL<643> A_IWL<642> A_IWL<641> A_IWL<640> A_IWL<639> A_IWL<638> A_IWL<637> A_IWL<636> A_IWL<635> A_IWL<634> A_IWL<633> A_IWL<632> A_IWL<631> A_IWL<630> A_IWL<629> A_IWL<628> A_IWL<627> A_IWL<626> A_IWL<625> A_IWL<624> A_IWL<623> A_IWL<622> A_IWL<621> A_IWL<620> A_IWL<619> A_IWL<618> A_IWL<617> A_IWL<616> A_IWL<615> A_IWL<614> A_IWL<613> A_IWL<612> A_IWL<611> A_IWL<610> A_IWL<609> A_IWL<608> A_IWL<607> A_IWL<606> A_IWL<605> A_IWL<604> A_IWL<603> A_IWL<602> A_IWL<601> A_IWL<600> A_IWL<599> A_IWL<598> A_IWL<597> A_IWL<596> A_IWL<595> A_IWL<594> A_IWL<593> A_IWL<592> A_IWL<591> A_IWL<590> A_IWL<589> A_IWL<588> A_IWL<587> A_IWL<586> A_IWL<585> A_IWL<584> A_IWL<583> A_IWL<582> A_IWL<581> A_IWL<580> A_IWL<579> A_IWL<578> A_IWL<577> A_IWL<576> A_IWL<575> A_IWL<574> A_IWL<573> A_IWL<572> A_IWL<571> A_IWL<570> A_IWL<569> A_IWL<568> A_IWL<567> A_IWL<566> A_IWL<565> A_IWL<564> A_IWL<563> A_IWL<562> A_IWL<561> A_IWL<560> A_IWL<559> A_IWL<558> A_IWL<557> A_IWL<556> A_IWL<555> A_IWL<554> A_IWL<553> A_IWL<552> A_IWL<551> A_IWL<550> A_IWL<549> A_IWL<548> A_IWL<547> A_IWL<546> A_IWL<545> A_IWL<544> A_IWL<543> A_IWL<542> A_IWL<541> A_IWL<540> A_IWL<539> A_IWL<538> A_IWL<537> A_IWL<536> A_IWL<535> A_IWL<534> A_IWL<533> A_IWL<532> A_IWL<531> A_IWL<530> A_IWL<529> A_IWL<528> A_IWL<527> A_IWL<526> A_IWL<525> A_IWL<524> A_IWL<523> A_IWL<522> A_IWL<521> A_IWL<520> A_IWL<519> A_IWL<518> A_IWL<517> A_IWL<516> A_IWL<515> A_IWL<514> A_IWL<513> A_IWL<512> A_IWL<1535> A_IWL<1534> A_IWL<1533> A_IWL<1532> A_IWL<1531> A_IWL<1530> A_IWL<1529> A_IWL<1528> A_IWL<1527> A_IWL<1526> A_IWL<1525> A_IWL<1524> A_IWL<1523> A_IWL<1522> A_IWL<1521> A_IWL<1520> A_IWL<1519> A_IWL<1518> A_IWL<1517> A_IWL<1516> A_IWL<1515> A_IWL<1514> A_IWL<1513> A_IWL<1512> A_IWL<1511> A_IWL<1510> A_IWL<1509> A_IWL<1508> A_IWL<1507> A_IWL<1506> A_IWL<1505> A_IWL<1504> A_IWL<1503> A_IWL<1502> A_IWL<1501> A_IWL<1500> A_IWL<1499> A_IWL<1498> A_IWL<1497> A_IWL<1496> A_IWL<1495> A_IWL<1494> A_IWL<1493> A_IWL<1492> A_IWL<1491> A_IWL<1490> A_IWL<1489> A_IWL<1488> A_IWL<1487> A_IWL<1486> A_IWL<1485> A_IWL<1484> A_IWL<1483> A_IWL<1482> A_IWL<1481> A_IWL<1480> A_IWL<1479> A_IWL<1478> A_IWL<1477> A_IWL<1476> A_IWL<1475> A_IWL<1474> A_IWL<1473> A_IWL<1472> A_IWL<1471> A_IWL<1470> A_IWL<1469> A_IWL<1468> A_IWL<1467> A_IWL<1466> A_IWL<1465> A_IWL<1464> A_IWL<1463> A_IWL<1462> A_IWL<1461> A_IWL<1460> A_IWL<1459> A_IWL<1458> A_IWL<1457> A_IWL<1456> A_IWL<1455> A_IWL<1454> A_IWL<1453> A_IWL<1452> A_IWL<1451> A_IWL<1450> A_IWL<1449> A_IWL<1448> A_IWL<1447> A_IWL<1446> A_IWL<1445> A_IWL<1444> A_IWL<1443> A_IWL<1442> A_IWL<1441> A_IWL<1440> A_IWL<1439> A_IWL<1438> A_IWL<1437> A_IWL<1436> A_IWL<1435> A_IWL<1434> A_IWL<1433> A_IWL<1432> A_IWL<1431> A_IWL<1430> A_IWL<1429> A_IWL<1428> A_IWL<1427> A_IWL<1426> A_IWL<1425> A_IWL<1424> A_IWL<1423> A_IWL<1422> A_IWL<1421> A_IWL<1420> A_IWL<1419> A_IWL<1418> A_IWL<1417> A_IWL<1416> A_IWL<1415> A_IWL<1414> A_IWL<1413> A_IWL<1412> A_IWL<1411> A_IWL<1410> A_IWL<1409> A_IWL<1408> A_IWL<1407> A_IWL<1406> A_IWL<1405> A_IWL<1404> A_IWL<1403> A_IWL<1402> A_IWL<1401> A_IWL<1400> A_IWL<1399> A_IWL<1398> A_IWL<1397> A_IWL<1396> A_IWL<1395> A_IWL<1394> A_IWL<1393> A_IWL<1392> A_IWL<1391> A_IWL<1390> A_IWL<1389> A_IWL<1388> A_IWL<1387> A_IWL<1386> A_IWL<1385> A_IWL<1384> A_IWL<1383> A_IWL<1382> A_IWL<1381> A_IWL<1380> A_IWL<1379> A_IWL<1378> A_IWL<1377> A_IWL<1376> A_IWL<1375> A_IWL<1374> A_IWL<1373> A_IWL<1372> A_IWL<1371> A_IWL<1370> A_IWL<1369> A_IWL<1368> A_IWL<1367> A_IWL<1366> A_IWL<1365> A_IWL<1364> A_IWL<1363> A_IWL<1362> A_IWL<1361> A_IWL<1360> A_IWL<1359> A_IWL<1358> A_IWL<1357> A_IWL<1356> A_IWL<1355> A_IWL<1354> A_IWL<1353> A_IWL<1352> A_IWL<1351> A_IWL<1350> A_IWL<1349> A_IWL<1348> A_IWL<1347> A_IWL<1346> A_IWL<1345> A_IWL<1344> A_IWL<1343> A_IWL<1342> A_IWL<1341> A_IWL<1340> A_IWL<1339> A_IWL<1338> A_IWL<1337> A_IWL<1336> A_IWL<1335> A_IWL<1334> A_IWL<1333> A_IWL<1332> A_IWL<1331> A_IWL<1330> A_IWL<1329> A_IWL<1328> A_IWL<1327> A_IWL<1326> A_IWL<1325> A_IWL<1324> A_IWL<1323> A_IWL<1322> A_IWL<1321> A_IWL<1320> A_IWL<1319> A_IWL<1318> A_IWL<1317> A_IWL<1316> A_IWL<1315> A_IWL<1314> A_IWL<1313> A_IWL<1312> A_IWL<1311> A_IWL<1310> A_IWL<1309> A_IWL<1308> A_IWL<1307> A_IWL<1306> A_IWL<1305> A_IWL<1304> A_IWL<1303> A_IWL<1302> A_IWL<1301> A_IWL<1300> A_IWL<1299> A_IWL<1298> A_IWL<1297> A_IWL<1296> A_IWL<1295> A_IWL<1294> A_IWL<1293> A_IWL<1292> A_IWL<1291> A_IWL<1290> A_IWL<1289> A_IWL<1288> A_IWL<1287> A_IWL<1286> A_IWL<1285> A_IWL<1284> A_IWL<1283> A_IWL<1282> A_IWL<1281> A_IWL<1280> A_IWL<1279> A_IWL<1278> A_IWL<1277> A_IWL<1276> A_IWL<1275> A_IWL<1274> A_IWL<1273> A_IWL<1272> A_IWL<1271> A_IWL<1270> A_IWL<1269> A_IWL<1268> A_IWL<1267> A_IWL<1266> A_IWL<1265> A_IWL<1264> A_IWL<1263> A_IWL<1262> A_IWL<1261> A_IWL<1260> A_IWL<1259> A_IWL<1258> A_IWL<1257> A_IWL<1256> A_IWL<1255> A_IWL<1254> A_IWL<1253> A_IWL<1252> A_IWL<1251> A_IWL<1250> A_IWL<1249> A_IWL<1248> A_IWL<1247> A_IWL<1246> A_IWL<1245> A_IWL<1244> A_IWL<1243> A_IWL<1242> A_IWL<1241> A_IWL<1240> A_IWL<1239> A_IWL<1238> A_IWL<1237> A_IWL<1236> A_IWL<1235> A_IWL<1234> A_IWL<1233> A_IWL<1232> A_IWL<1231> A_IWL<1230> A_IWL<1229> A_IWL<1228> A_IWL<1227> A_IWL<1226> A_IWL<1225> A_IWL<1224> A_IWL<1223> A_IWL<1222> A_IWL<1221> A_IWL<1220> A_IWL<1219> A_IWL<1218> A_IWL<1217> A_IWL<1216> A_IWL<1215> A_IWL<1214> A_IWL<1213> A_IWL<1212> A_IWL<1211> A_IWL<1210> A_IWL<1209> A_IWL<1208> A_IWL<1207> A_IWL<1206> A_IWL<1205> A_IWL<1204> A_IWL<1203> A_IWL<1202> A_IWL<1201> A_IWL<1200> A_IWL<1199> A_IWL<1198> A_IWL<1197> A_IWL<1196> A_IWL<1195> A_IWL<1194> A_IWL<1193> A_IWL<1192> A_IWL<1191> A_IWL<1190> A_IWL<1189> A_IWL<1188> A_IWL<1187> A_IWL<1186> A_IWL<1185> A_IWL<1184> A_IWL<1183> A_IWL<1182> A_IWL<1181> A_IWL<1180> A_IWL<1179> A_IWL<1178> A_IWL<1177> A_IWL<1176> A_IWL<1175> A_IWL<1174> A_IWL<1173> A_IWL<1172> A_IWL<1171> A_IWL<1170> A_IWL<1169> A_IWL<1168> A_IWL<1167> A_IWL<1166> A_IWL<1165> A_IWL<1164> A_IWL<1163> A_IWL<1162> A_IWL<1161> A_IWL<1160> A_IWL<1159> A_IWL<1158> A_IWL<1157> A_IWL<1156> A_IWL<1155> A_IWL<1154> A_IWL<1153> A_IWL<1152> A_IWL<1151> A_IWL<1150> A_IWL<1149> A_IWL<1148> A_IWL<1147> A_IWL<1146> A_IWL<1145> A_IWL<1144> A_IWL<1143> A_IWL<1142> A_IWL<1141> A_IWL<1140> A_IWL<1139> A_IWL<1138> A_IWL<1137> A_IWL<1136> A_IWL<1135> A_IWL<1134> A_IWL<1133> A_IWL<1132> A_IWL<1131> A_IWL<1130> A_IWL<1129> A_IWL<1128> A_IWL<1127> A_IWL<1126> A_IWL<1125> A_IWL<1124> A_IWL<1123> A_IWL<1122> A_IWL<1121> A_IWL<1120> A_IWL<1119> A_IWL<1118> A_IWL<1117> A_IWL<1116> A_IWL<1115> A_IWL<1114> A_IWL<1113> A_IWL<1112> A_IWL<1111> A_IWL<1110> A_IWL<1109> A_IWL<1108> A_IWL<1107> A_IWL<1106> A_IWL<1105> A_IWL<1104> A_IWL<1103> A_IWL<1102> A_IWL<1101> A_IWL<1100> A_IWL<1099> A_IWL<1098> A_IWL<1097> A_IWL<1096> A_IWL<1095> A_IWL<1094> A_IWL<1093> A_IWL<1092> A_IWL<1091> A_IWL<1090> A_IWL<1089> A_IWL<1088> A_IWL<1087> A_IWL<1086> A_IWL<1085> A_IWL<1084> A_IWL<1083> A_IWL<1082> A_IWL<1081> A_IWL<1080> A_IWL<1079> A_IWL<1078> A_IWL<1077> A_IWL<1076> A_IWL<1075> A_IWL<1074> A_IWL<1073> A_IWL<1072> A_IWL<1071> A_IWL<1070> A_IWL<1069> A_IWL<1068> A_IWL<1067> A_IWL<1066> A_IWL<1065> A_IWL<1064> A_IWL<1063> A_IWL<1062> A_IWL<1061> A_IWL<1060> A_IWL<1059> A_IWL<1058> A_IWL<1057> A_IWL<1056> A_IWL<1055> A_IWL<1054> A_IWL<1053> A_IWL<1052> A_IWL<1051> A_IWL<1050> A_IWL<1049> A_IWL<1048> A_IWL<1047> A_IWL<1046> A_IWL<1045> A_IWL<1044> A_IWL<1043> A_IWL<1042> A_IWL<1041> A_IWL<1040> A_IWL<1039> A_IWL<1038> A_IWL<1037> A_IWL<1036> A_IWL<1035> A_IWL<1034> A_IWL<1033> A_IWL<1032> A_IWL<1031> A_IWL<1030> A_IWL<1029> A_IWL<1028> A_IWL<1027> A_IWL<1026> A_IWL<1025> A_IWL<1024> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<1> A_BLC<3> A_BLC<2> A_BLC_TOP<3> A_BLC_TOP<2> A_BLT<3> A_BLT<2> A_BLT_TOP<3> A_BLT_TOP<2> A_IWL<511> A_IWL<510> A_IWL<509> A_IWL<508> A_IWL<507> A_IWL<506> A_IWL<505> A_IWL<504> A_IWL<503> A_IWL<502> A_IWL<501> A_IWL<500> A_IWL<499> A_IWL<498> A_IWL<497> A_IWL<496> A_IWL<495> A_IWL<494> A_IWL<493> A_IWL<492> A_IWL<491> A_IWL<490> A_IWL<489> A_IWL<488> A_IWL<487> A_IWL<486> A_IWL<485> A_IWL<484> A_IWL<483> A_IWL<482> A_IWL<481> A_IWL<480> A_IWL<479> A_IWL<478> A_IWL<477> A_IWL<476> A_IWL<475> A_IWL<474> A_IWL<473> A_IWL<472> A_IWL<471> A_IWL<470> A_IWL<469> A_IWL<468> A_IWL<467> A_IWL<466> A_IWL<465> A_IWL<464> A_IWL<463> A_IWL<462> A_IWL<461> A_IWL<460> A_IWL<459> A_IWL<458> A_IWL<457> A_IWL<456> A_IWL<455> A_IWL<454> A_IWL<453> A_IWL<452> A_IWL<451> A_IWL<450> A_IWL<449> A_IWL<448> A_IWL<447> A_IWL<446> A_IWL<445> A_IWL<444> A_IWL<443> A_IWL<442> A_IWL<441> A_IWL<440> A_IWL<439> A_IWL<438> A_IWL<437> A_IWL<436> A_IWL<435> A_IWL<434> A_IWL<433> A_IWL<432> A_IWL<431> A_IWL<430> A_IWL<429> A_IWL<428> A_IWL<427> A_IWL<426> A_IWL<425> A_IWL<424> A_IWL<423> A_IWL<422> A_IWL<421> A_IWL<420> A_IWL<419> A_IWL<418> A_IWL<417> A_IWL<416> A_IWL<415> A_IWL<414> A_IWL<413> A_IWL<412> A_IWL<411> A_IWL<410> A_IWL<409> A_IWL<408> A_IWL<407> A_IWL<406> A_IWL<405> A_IWL<404> A_IWL<403> A_IWL<402> A_IWL<401> A_IWL<400> A_IWL<399> A_IWL<398> A_IWL<397> A_IWL<396> A_IWL<395> A_IWL<394> A_IWL<393> A_IWL<392> A_IWL<391> A_IWL<390> A_IWL<389> A_IWL<388> A_IWL<387> A_IWL<386> A_IWL<385> A_IWL<384> A_IWL<383> A_IWL<382> A_IWL<381> A_IWL<380> A_IWL<379> A_IWL<378> A_IWL<377> A_IWL<376> A_IWL<375> A_IWL<374> A_IWL<373> A_IWL<372> A_IWL<371> A_IWL<370> A_IWL<369> A_IWL<368> A_IWL<367> A_IWL<366> A_IWL<365> A_IWL<364> A_IWL<363> A_IWL<362> A_IWL<361> A_IWL<360> A_IWL<359> A_IWL<358> A_IWL<357> A_IWL<356> A_IWL<355> A_IWL<354> A_IWL<353> A_IWL<352> A_IWL<351> A_IWL<350> A_IWL<349> A_IWL<348> A_IWL<347> A_IWL<346> A_IWL<345> A_IWL<344> A_IWL<343> A_IWL<342> A_IWL<341> A_IWL<340> A_IWL<339> A_IWL<338> A_IWL<337> A_IWL<336> A_IWL<335> A_IWL<334> A_IWL<333> A_IWL<332> A_IWL<331> A_IWL<330> A_IWL<329> A_IWL<328> A_IWL<327> A_IWL<326> A_IWL<325> A_IWL<324> A_IWL<323> A_IWL<322> A_IWL<321> A_IWL<320> A_IWL<319> A_IWL<318> A_IWL<317> A_IWL<316> A_IWL<315> A_IWL<314> A_IWL<313> A_IWL<312> A_IWL<311> A_IWL<310> A_IWL<309> A_IWL<308> A_IWL<307> A_IWL<306> A_IWL<305> A_IWL<304> A_IWL<303> A_IWL<302> A_IWL<301> A_IWL<300> A_IWL<299> A_IWL<298> A_IWL<297> A_IWL<296> A_IWL<295> A_IWL<294> A_IWL<293> A_IWL<292> A_IWL<291> A_IWL<290> A_IWL<289> A_IWL<288> A_IWL<287> A_IWL<286> A_IWL<285> A_IWL<284> A_IWL<283> A_IWL<282> A_IWL<281> A_IWL<280> A_IWL<279> A_IWL<278> A_IWL<277> A_IWL<276> A_IWL<275> A_IWL<274> A_IWL<273> A_IWL<272> A_IWL<271> A_IWL<270> A_IWL<269> A_IWL<268> A_IWL<267> A_IWL<266> A_IWL<265> A_IWL<264> A_IWL<263> A_IWL<262> A_IWL<261> A_IWL<260> A_IWL<259> A_IWL<258> A_IWL<257> A_IWL<256> A_IWL<255> A_IWL<254> A_IWL<253> A_IWL<252> A_IWL<251> A_IWL<250> A_IWL<249> A_IWL<248> A_IWL<247> A_IWL<246> A_IWL<245> A_IWL<244> A_IWL<243> A_IWL<242> A_IWL<241> A_IWL<240> A_IWL<239> A_IWL<238> A_IWL<237> A_IWL<236> A_IWL<235> A_IWL<234> A_IWL<233> A_IWL<232> A_IWL<231> A_IWL<230> A_IWL<229> A_IWL<228> A_IWL<227> A_IWL<226> A_IWL<225> A_IWL<224> A_IWL<223> A_IWL<222> A_IWL<221> A_IWL<220> A_IWL<219> A_IWL<218> A_IWL<217> A_IWL<216> A_IWL<215> A_IWL<214> A_IWL<213> A_IWL<212> A_IWL<211> A_IWL<210> A_IWL<209> A_IWL<208> A_IWL<207> A_IWL<206> A_IWL<205> A_IWL<204> A_IWL<203> A_IWL<202> A_IWL<201> A_IWL<200> A_IWL<199> A_IWL<198> A_IWL<197> A_IWL<196> A_IWL<195> A_IWL<194> A_IWL<193> A_IWL<192> A_IWL<191> A_IWL<190> A_IWL<189> A_IWL<188> A_IWL<187> A_IWL<186> A_IWL<185> A_IWL<184> A_IWL<183> A_IWL<182> A_IWL<181> A_IWL<180> A_IWL<179> A_IWL<178> A_IWL<177> A_IWL<176> A_IWL<175> A_IWL<174> A_IWL<173> A_IWL<172> A_IWL<171> A_IWL<170> A_IWL<169> A_IWL<168> A_IWL<167> A_IWL<166> A_IWL<165> A_IWL<164> A_IWL<163> A_IWL<162> A_IWL<161> A_IWL<160> A_IWL<159> A_IWL<158> A_IWL<157> A_IWL<156> A_IWL<155> A_IWL<154> A_IWL<153> A_IWL<152> A_IWL<151> A_IWL<150> A_IWL<149> A_IWL<148> A_IWL<147> A_IWL<146> A_IWL<145> A_IWL<144> A_IWL<143> A_IWL<142> A_IWL<141> A_IWL<140> A_IWL<139> A_IWL<138> A_IWL<137> A_IWL<136> A_IWL<135> A_IWL<134> A_IWL<133> A_IWL<132> A_IWL<131> A_IWL<130> A_IWL<129> A_IWL<128> A_IWL<127> A_IWL<126> A_IWL<125> A_IWL<124> A_IWL<123> A_IWL<122> A_IWL<121> A_IWL<120> A_IWL<119> A_IWL<118> A_IWL<117> A_IWL<116> A_IWL<115> A_IWL<114> A_IWL<113> A_IWL<112> A_IWL<111> A_IWL<110> A_IWL<109> A_IWL<108> A_IWL<107> A_IWL<106> A_IWL<105> A_IWL<104> A_IWL<103> A_IWL<102> A_IWL<101> A_IWL<100> A_IWL<99> A_IWL<98> A_IWL<97> A_IWL<96> A_IWL<95> A_IWL<94> A_IWL<93> A_IWL<92> A_IWL<91> A_IWL<90> A_IWL<89> A_IWL<88> A_IWL<87> A_IWL<86> A_IWL<85> A_IWL<84> A_IWL<83> A_IWL<82> A_IWL<81> A_IWL<80> A_IWL<79> A_IWL<78> A_IWL<77> A_IWL<76> A_IWL<75> A_IWL<74> A_IWL<73> A_IWL<72> A_IWL<71> A_IWL<70> A_IWL<69> A_IWL<68> A_IWL<67> A_IWL<66> A_IWL<65> A_IWL<64> A_IWL<63> A_IWL<62> A_IWL<61> A_IWL<60> A_IWL<59> A_IWL<58> A_IWL<57> A_IWL<56> A_IWL<55> A_IWL<54> A_IWL<53> A_IWL<52> A_IWL<51> A_IWL<50> A_IWL<49> A_IWL<48> A_IWL<47> A_IWL<46> A_IWL<45> A_IWL<44> A_IWL<43> A_IWL<42> A_IWL<41> A_IWL<40> A_IWL<39> A_IWL<38> A_IWL<37> A_IWL<36> A_IWL<35> A_IWL<34> A_IWL<33> A_IWL<32> A_IWL<31> A_IWL<30> A_IWL<29> A_IWL<28> A_IWL<27> A_IWL<26> A_IWL<25> A_IWL<24> A_IWL<23> A_IWL<22> A_IWL<21> A_IWL<20> A_IWL<19> A_IWL<18> A_IWL<17> A_IWL<16> A_IWL<15> A_IWL<14> A_IWL<13> A_IWL<12> A_IWL<11> A_IWL<10> A_IWL<9> A_IWL<8> A_IWL<7> A_IWL<6> A_IWL<5> A_IWL<4> A_IWL<3> A_IWL<2> A_IWL<1> A_IWL<0> A_IWL<1023> A_IWL<1022> A_IWL<1021> A_IWL<1020> A_IWL<1019> A_IWL<1018> A_IWL<1017> A_IWL<1016> A_IWL<1015> A_IWL<1014> A_IWL<1013> A_IWL<1012> A_IWL<1011> A_IWL<1010> A_IWL<1009> A_IWL<1008> A_IWL<1007> A_IWL<1006> A_IWL<1005> A_IWL<1004> A_IWL<1003> A_IWL<1002> A_IWL<1001> A_IWL<1000> A_IWL<999> A_IWL<998> A_IWL<997> A_IWL<996> A_IWL<995> A_IWL<994> A_IWL<993> A_IWL<992> A_IWL<991> A_IWL<990> A_IWL<989> A_IWL<988> A_IWL<987> A_IWL<986> A_IWL<985> A_IWL<984> A_IWL<983> A_IWL<982> A_IWL<981> A_IWL<980> A_IWL<979> A_IWL<978> A_IWL<977> A_IWL<976> A_IWL<975> A_IWL<974> A_IWL<973> A_IWL<972> A_IWL<971> A_IWL<970> A_IWL<969> A_IWL<968> A_IWL<967> A_IWL<966> A_IWL<965> A_IWL<964> A_IWL<963> A_IWL<962> A_IWL<961> A_IWL<960> A_IWL<959> A_IWL<958> A_IWL<957> A_IWL<956> A_IWL<955> A_IWL<954> A_IWL<953> A_IWL<952> A_IWL<951> A_IWL<950> A_IWL<949> A_IWL<948> A_IWL<947> A_IWL<946> A_IWL<945> A_IWL<944> A_IWL<943> A_IWL<942> A_IWL<941> A_IWL<940> A_IWL<939> A_IWL<938> A_IWL<937> A_IWL<936> A_IWL<935> A_IWL<934> A_IWL<933> A_IWL<932> A_IWL<931> A_IWL<930> A_IWL<929> A_IWL<928> A_IWL<927> A_IWL<926> A_IWL<925> A_IWL<924> A_IWL<923> A_IWL<922> A_IWL<921> A_IWL<920> A_IWL<919> A_IWL<918> A_IWL<917> A_IWL<916> A_IWL<915> A_IWL<914> A_IWL<913> A_IWL<912> A_IWL<911> A_IWL<910> A_IWL<909> A_IWL<908> A_IWL<907> A_IWL<906> A_IWL<905> A_IWL<904> A_IWL<903> A_IWL<902> A_IWL<901> A_IWL<900> A_IWL<899> A_IWL<898> A_IWL<897> A_IWL<896> A_IWL<895> A_IWL<894> A_IWL<893> A_IWL<892> A_IWL<891> A_IWL<890> A_IWL<889> A_IWL<888> A_IWL<887> A_IWL<886> A_IWL<885> A_IWL<884> A_IWL<883> A_IWL<882> A_IWL<881> A_IWL<880> A_IWL<879> A_IWL<878> A_IWL<877> A_IWL<876> A_IWL<875> A_IWL<874> A_IWL<873> A_IWL<872> A_IWL<871> A_IWL<870> A_IWL<869> A_IWL<868> A_IWL<867> A_IWL<866> A_IWL<865> A_IWL<864> A_IWL<863> A_IWL<862> A_IWL<861> A_IWL<860> A_IWL<859> A_IWL<858> A_IWL<857> A_IWL<856> A_IWL<855> A_IWL<854> A_IWL<853> A_IWL<852> A_IWL<851> A_IWL<850> A_IWL<849> A_IWL<848> A_IWL<847> A_IWL<846> A_IWL<845> A_IWL<844> A_IWL<843> A_IWL<842> A_IWL<841> A_IWL<840> A_IWL<839> A_IWL<838> A_IWL<837> A_IWL<836> A_IWL<835> A_IWL<834> A_IWL<833> A_IWL<832> A_IWL<831> A_IWL<830> A_IWL<829> A_IWL<828> A_IWL<827> A_IWL<826> A_IWL<825> A_IWL<824> A_IWL<823> A_IWL<822> A_IWL<821> A_IWL<820> A_IWL<819> A_IWL<818> A_IWL<817> A_IWL<816> A_IWL<815> A_IWL<814> A_IWL<813> A_IWL<812> A_IWL<811> A_IWL<810> A_IWL<809> A_IWL<808> A_IWL<807> A_IWL<806> A_IWL<805> A_IWL<804> A_IWL<803> A_IWL<802> A_IWL<801> A_IWL<800> A_IWL<799> A_IWL<798> A_IWL<797> A_IWL<796> A_IWL<795> A_IWL<794> A_IWL<793> A_IWL<792> A_IWL<791> A_IWL<790> A_IWL<789> A_IWL<788> A_IWL<787> A_IWL<786> A_IWL<785> A_IWL<784> A_IWL<783> A_IWL<782> A_IWL<781> A_IWL<780> A_IWL<779> A_IWL<778> A_IWL<777> A_IWL<776> A_IWL<775> A_IWL<774> A_IWL<773> A_IWL<772> A_IWL<771> A_IWL<770> A_IWL<769> A_IWL<768> A_IWL<767> A_IWL<766> A_IWL<765> A_IWL<764> A_IWL<763> A_IWL<762> A_IWL<761> A_IWL<760> A_IWL<759> A_IWL<758> A_IWL<757> A_IWL<756> A_IWL<755> A_IWL<754> A_IWL<753> A_IWL<752> A_IWL<751> A_IWL<750> A_IWL<749> A_IWL<748> A_IWL<747> A_IWL<746> A_IWL<745> A_IWL<744> A_IWL<743> A_IWL<742> A_IWL<741> A_IWL<740> A_IWL<739> A_IWL<738> A_IWL<737> A_IWL<736> A_IWL<735> A_IWL<734> A_IWL<733> A_IWL<732> A_IWL<731> A_IWL<730> A_IWL<729> A_IWL<728> A_IWL<727> A_IWL<726> A_IWL<725> A_IWL<724> A_IWL<723> A_IWL<722> A_IWL<721> A_IWL<720> A_IWL<719> A_IWL<718> A_IWL<717> A_IWL<716> A_IWL<715> A_IWL<714> A_IWL<713> A_IWL<712> A_IWL<711> A_IWL<710> A_IWL<709> A_IWL<708> A_IWL<707> A_IWL<706> A_IWL<705> A_IWL<704> A_IWL<703> A_IWL<702> A_IWL<701> A_IWL<700> A_IWL<699> A_IWL<698> A_IWL<697> A_IWL<696> A_IWL<695> A_IWL<694> A_IWL<693> A_IWL<692> A_IWL<691> A_IWL<690> A_IWL<689> A_IWL<688> A_IWL<687> A_IWL<686> A_IWL<685> A_IWL<684> A_IWL<683> A_IWL<682> A_IWL<681> A_IWL<680> A_IWL<679> A_IWL<678> A_IWL<677> A_IWL<676> A_IWL<675> A_IWL<674> A_IWL<673> A_IWL<672> A_IWL<671> A_IWL<670> A_IWL<669> A_IWL<668> A_IWL<667> A_IWL<666> A_IWL<665> A_IWL<664> A_IWL<663> A_IWL<662> A_IWL<661> A_IWL<660> A_IWL<659> A_IWL<658> A_IWL<657> A_IWL<656> A_IWL<655> A_IWL<654> A_IWL<653> A_IWL<652> A_IWL<651> A_IWL<650> A_IWL<649> A_IWL<648> A_IWL<647> A_IWL<646> A_IWL<645> A_IWL<644> A_IWL<643> A_IWL<642> A_IWL<641> A_IWL<640> A_IWL<639> A_IWL<638> A_IWL<637> A_IWL<636> A_IWL<635> A_IWL<634> A_IWL<633> A_IWL<632> A_IWL<631> A_IWL<630> A_IWL<629> A_IWL<628> A_IWL<627> A_IWL<626> A_IWL<625> A_IWL<624> A_IWL<623> A_IWL<622> A_IWL<621> A_IWL<620> A_IWL<619> A_IWL<618> A_IWL<617> A_IWL<616> A_IWL<615> A_IWL<614> A_IWL<613> A_IWL<612> A_IWL<611> A_IWL<610> A_IWL<609> A_IWL<608> A_IWL<607> A_IWL<606> A_IWL<605> A_IWL<604> A_IWL<603> A_IWL<602> A_IWL<601> A_IWL<600> A_IWL<599> A_IWL<598> A_IWL<597> A_IWL<596> A_IWL<595> A_IWL<594> A_IWL<593> A_IWL<592> A_IWL<591> A_IWL<590> A_IWL<589> A_IWL<588> A_IWL<587> A_IWL<586> A_IWL<585> A_IWL<584> A_IWL<583> A_IWL<582> A_IWL<581> A_IWL<580> A_IWL<579> A_IWL<578> A_IWL<577> A_IWL<576> A_IWL<575> A_IWL<574> A_IWL<573> A_IWL<572> A_IWL<571> A_IWL<570> A_IWL<569> A_IWL<568> A_IWL<567> A_IWL<566> A_IWL<565> A_IWL<564> A_IWL<563> A_IWL<562> A_IWL<561> A_IWL<560> A_IWL<559> A_IWL<558> A_IWL<557> A_IWL<556> A_IWL<555> A_IWL<554> A_IWL<553> A_IWL<552> A_IWL<551> A_IWL<550> A_IWL<549> A_IWL<548> A_IWL<547> A_IWL<546> A_IWL<545> A_IWL<544> A_IWL<543> A_IWL<542> A_IWL<541> A_IWL<540> A_IWL<539> A_IWL<538> A_IWL<537> A_IWL<536> A_IWL<535> A_IWL<534> A_IWL<533> A_IWL<532> A_IWL<531> A_IWL<530> A_IWL<529> A_IWL<528> A_IWL<527> A_IWL<526> A_IWL<525> A_IWL<524> A_IWL<523> A_IWL<522> A_IWL<521> A_IWL<520> A_IWL<519> A_IWL<518> A_IWL<517> A_IWL<516> A_IWL<515> A_IWL<514> A_IWL<513> A_IWL<512> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
XCOL<0> A_BLC<1> A_BLC<0> A_BLC_TOP<1> A_BLC_TOP<0> A_BLT<1> A_BLT<0> A_BLT_TOP<1> A_BLT_TOP<0> A_WL<511> A_WL<510> A_WL<509> A_WL<508> A_WL<507> A_WL<506> A_WL<505> A_WL<504> A_WL<503> A_WL<502> A_WL<501> A_WL<500> A_WL<499> A_WL<498> A_WL<497> A_WL<496> A_WL<495> A_WL<494> A_WL<493> A_WL<492> A_WL<491> A_WL<490> A_WL<489> A_WL<488> A_WL<487> A_WL<486> A_WL<485> A_WL<484> A_WL<483> A_WL<482> A_WL<481> A_WL<480> A_WL<479> A_WL<478> A_WL<477> A_WL<476> A_WL<475> A_WL<474> A_WL<473> A_WL<472> A_WL<471> A_WL<470> A_WL<469> A_WL<468> A_WL<467> A_WL<466> A_WL<465> A_WL<464> A_WL<463> A_WL<462> A_WL<461> A_WL<460> A_WL<459> A_WL<458> A_WL<457> A_WL<456> A_WL<455> A_WL<454> A_WL<453> A_WL<452> A_WL<451> A_WL<450> A_WL<449> A_WL<448> A_WL<447> A_WL<446> A_WL<445> A_WL<444> A_WL<443> A_WL<442> A_WL<441> A_WL<440> A_WL<439> A_WL<438> A_WL<437> A_WL<436> A_WL<435> A_WL<434> A_WL<433> A_WL<432> A_WL<431> A_WL<430> A_WL<429> A_WL<428> A_WL<427> A_WL<426> A_WL<425> A_WL<424> A_WL<423> A_WL<422> A_WL<421> A_WL<420> A_WL<419> A_WL<418> A_WL<417> A_WL<416> A_WL<415> A_WL<414> A_WL<413> A_WL<412> A_WL<411> A_WL<410> A_WL<409> A_WL<408> A_WL<407> A_WL<406> A_WL<405> A_WL<404> A_WL<403> A_WL<402> A_WL<401> A_WL<400> A_WL<399> A_WL<398> A_WL<397> A_WL<396> A_WL<395> A_WL<394> A_WL<393> A_WL<392> A_WL<391> A_WL<390> A_WL<389> A_WL<388> A_WL<387> A_WL<386> A_WL<385> A_WL<384> A_WL<383> A_WL<382> A_WL<381> A_WL<380> A_WL<379> A_WL<378> A_WL<377> A_WL<376> A_WL<375> A_WL<374> A_WL<373> A_WL<372> A_WL<371> A_WL<370> A_WL<369> A_WL<368> A_WL<367> A_WL<366> A_WL<365> A_WL<364> A_WL<363> A_WL<362> A_WL<361> A_WL<360> A_WL<359> A_WL<358> A_WL<357> A_WL<356> A_WL<355> A_WL<354> A_WL<353> A_WL<352> A_WL<351> A_WL<350> A_WL<349> A_WL<348> A_WL<347> A_WL<346> A_WL<345> A_WL<344> A_WL<343> A_WL<342> A_WL<341> A_WL<340> A_WL<339> A_WL<338> A_WL<337> A_WL<336> A_WL<335> A_WL<334> A_WL<333> A_WL<332> A_WL<331> A_WL<330> A_WL<329> A_WL<328> A_WL<327> A_WL<326> A_WL<325> A_WL<324> A_WL<323> A_WL<322> A_WL<321> A_WL<320> A_WL<319> A_WL<318> A_WL<317> A_WL<316> A_WL<315> A_WL<314> A_WL<313> A_WL<312> A_WL<311> A_WL<310> A_WL<309> A_WL<308> A_WL<307> A_WL<306> A_WL<305> A_WL<304> A_WL<303> A_WL<302> A_WL<301> A_WL<300> A_WL<299> A_WL<298> A_WL<297> A_WL<296> A_WL<295> A_WL<294> A_WL<293> A_WL<292> A_WL<291> A_WL<290> A_WL<289> A_WL<288> A_WL<287> A_WL<286> A_WL<285> A_WL<284> A_WL<283> A_WL<282> A_WL<281> A_WL<280> A_WL<279> A_WL<278> A_WL<277> A_WL<276> A_WL<275> A_WL<274> A_WL<273> A_WL<272> A_WL<271> A_WL<270> A_WL<269> A_WL<268> A_WL<267> A_WL<266> A_WL<265> A_WL<264> A_WL<263> A_WL<262> A_WL<261> A_WL<260> A_WL<259> A_WL<258> A_WL<257> A_WL<256> A_WL<255> A_WL<254> A_WL<253> A_WL<252> A_WL<251> A_WL<250> A_WL<249> A_WL<248> A_WL<247> A_WL<246> A_WL<245> A_WL<244> A_WL<243> A_WL<242> A_WL<241> A_WL<240> A_WL<239> A_WL<238> A_WL<237> A_WL<236> A_WL<235> A_WL<234> A_WL<233> A_WL<232> A_WL<231> A_WL<230> A_WL<229> A_WL<228> A_WL<227> A_WL<226> A_WL<225> A_WL<224> A_WL<223> A_WL<222> A_WL<221> A_WL<220> A_WL<219> A_WL<218> A_WL<217> A_WL<216> A_WL<215> A_WL<214> A_WL<213> A_WL<212> A_WL<211> A_WL<210> A_WL<209> A_WL<208> A_WL<207> A_WL<206> A_WL<205> A_WL<204> A_WL<203> A_WL<202> A_WL<201> A_WL<200> A_WL<199> A_WL<198> A_WL<197> A_WL<196> A_WL<195> A_WL<194> A_WL<193> A_WL<192> A_WL<191> A_WL<190> A_WL<189> A_WL<188> A_WL<187> A_WL<186> A_WL<185> A_WL<184> A_WL<183> A_WL<182> A_WL<181> A_WL<180> A_WL<179> A_WL<178> A_WL<177> A_WL<176> A_WL<175> A_WL<174> A_WL<173> A_WL<172> A_WL<171> A_WL<170> A_WL<169> A_WL<168> A_WL<167> A_WL<166> A_WL<165> A_WL<164> A_WL<163> A_WL<162> A_WL<161> A_WL<160> A_WL<159> A_WL<158> A_WL<157> A_WL<156> A_WL<155> A_WL<154> A_WL<153> A_WL<152> A_WL<151> A_WL<150> A_WL<149> A_WL<148> A_WL<147> A_WL<146> A_WL<145> A_WL<144> A_WL<143> A_WL<142> A_WL<141> A_WL<140> A_WL<139> A_WL<138> A_WL<137> A_WL<136> A_WL<135> A_WL<134> A_WL<133> A_WL<132> A_WL<131> A_WL<130> A_WL<129> A_WL<128> A_WL<127> A_WL<126> A_WL<125> A_WL<124> A_WL<123> A_WL<122> A_WL<121> A_WL<120> A_WL<119> A_WL<118> A_WL<117> A_WL<116> A_WL<115> A_WL<114> A_WL<113> A_WL<112> A_WL<111> A_WL<110> A_WL<109> A_WL<108> A_WL<107> A_WL<106> A_WL<105> A_WL<104> A_WL<103> A_WL<102> A_WL<101> A_WL<100> A_WL<99> A_WL<98> A_WL<97> A_WL<96> A_WL<95> A_WL<94> A_WL<93> A_WL<92> A_WL<91> A_WL<90> A_WL<89> A_WL<88> A_WL<87> A_WL<86> A_WL<85> A_WL<84> A_WL<83> A_WL<82> A_WL<81> A_WL<80> A_WL<79> A_WL<78> A_WL<77> A_WL<76> A_WL<75> A_WL<74> A_WL<73> A_WL<72> A_WL<71> A_WL<70> A_WL<69> A_WL<68> A_WL<67> A_WL<66> A_WL<65> A_WL<64> A_WL<63> A_WL<62> A_WL<61> A_WL<60> A_WL<59> A_WL<58> A_WL<57> A_WL<56> A_WL<55> A_WL<54> A_WL<53> A_WL<52> A_WL<51> A_WL<50> A_WL<49> A_WL<48> A_WL<47> A_WL<46> A_WL<45> A_WL<44> A_WL<43> A_WL<42> A_WL<41> A_WL<40> A_WL<39> A_WL<38> A_WL<37> A_WL<36> A_WL<35> A_WL<34> A_WL<33> A_WL<32> A_WL<31> A_WL<30> A_WL<29> A_WL<28> A_WL<27> A_WL<26> A_WL<25> A_WL<24> A_WL<23> A_WL<22> A_WL<21> A_WL<20> A_WL<19> A_WL<18> A_WL<17> A_WL<16> A_WL<15> A_WL<14> A_WL<13> A_WL<12> A_WL<11> A_WL<10> A_WL<9> A_WL<8> A_WL<7> A_WL<6> A_WL<5> A_WL<4> A_WL<3> A_WL<2> A_WL<1> A_WL<0> A_IWL<511> A_IWL<510> A_IWL<509> A_IWL<508> A_IWL<507> A_IWL<506> A_IWL<505> A_IWL<504> A_IWL<503> A_IWL<502> A_IWL<501> A_IWL<500> A_IWL<499> A_IWL<498> A_IWL<497> A_IWL<496> A_IWL<495> A_IWL<494> A_IWL<493> A_IWL<492> A_IWL<491> A_IWL<490> A_IWL<489> A_IWL<488> A_IWL<487> A_IWL<486> A_IWL<485> A_IWL<484> A_IWL<483> A_IWL<482> A_IWL<481> A_IWL<480> A_IWL<479> A_IWL<478> A_IWL<477> A_IWL<476> A_IWL<475> A_IWL<474> A_IWL<473> A_IWL<472> A_IWL<471> A_IWL<470> A_IWL<469> A_IWL<468> A_IWL<467> A_IWL<466> A_IWL<465> A_IWL<464> A_IWL<463> A_IWL<462> A_IWL<461> A_IWL<460> A_IWL<459> A_IWL<458> A_IWL<457> A_IWL<456> A_IWL<455> A_IWL<454> A_IWL<453> A_IWL<452> A_IWL<451> A_IWL<450> A_IWL<449> A_IWL<448> A_IWL<447> A_IWL<446> A_IWL<445> A_IWL<444> A_IWL<443> A_IWL<442> A_IWL<441> A_IWL<440> A_IWL<439> A_IWL<438> A_IWL<437> A_IWL<436> A_IWL<435> A_IWL<434> A_IWL<433> A_IWL<432> A_IWL<431> A_IWL<430> A_IWL<429> A_IWL<428> A_IWL<427> A_IWL<426> A_IWL<425> A_IWL<424> A_IWL<423> A_IWL<422> A_IWL<421> A_IWL<420> A_IWL<419> A_IWL<418> A_IWL<417> A_IWL<416> A_IWL<415> A_IWL<414> A_IWL<413> A_IWL<412> A_IWL<411> A_IWL<410> A_IWL<409> A_IWL<408> A_IWL<407> A_IWL<406> A_IWL<405> A_IWL<404> A_IWL<403> A_IWL<402> A_IWL<401> A_IWL<400> A_IWL<399> A_IWL<398> A_IWL<397> A_IWL<396> A_IWL<395> A_IWL<394> A_IWL<393> A_IWL<392> A_IWL<391> A_IWL<390> A_IWL<389> A_IWL<388> A_IWL<387> A_IWL<386> A_IWL<385> A_IWL<384> A_IWL<383> A_IWL<382> A_IWL<381> A_IWL<380> A_IWL<379> A_IWL<378> A_IWL<377> A_IWL<376> A_IWL<375> A_IWL<374> A_IWL<373> A_IWL<372> A_IWL<371> A_IWL<370> A_IWL<369> A_IWL<368> A_IWL<367> A_IWL<366> A_IWL<365> A_IWL<364> A_IWL<363> A_IWL<362> A_IWL<361> A_IWL<360> A_IWL<359> A_IWL<358> A_IWL<357> A_IWL<356> A_IWL<355> A_IWL<354> A_IWL<353> A_IWL<352> A_IWL<351> A_IWL<350> A_IWL<349> A_IWL<348> A_IWL<347> A_IWL<346> A_IWL<345> A_IWL<344> A_IWL<343> A_IWL<342> A_IWL<341> A_IWL<340> A_IWL<339> A_IWL<338> A_IWL<337> A_IWL<336> A_IWL<335> A_IWL<334> A_IWL<333> A_IWL<332> A_IWL<331> A_IWL<330> A_IWL<329> A_IWL<328> A_IWL<327> A_IWL<326> A_IWL<325> A_IWL<324> A_IWL<323> A_IWL<322> A_IWL<321> A_IWL<320> A_IWL<319> A_IWL<318> A_IWL<317> A_IWL<316> A_IWL<315> A_IWL<314> A_IWL<313> A_IWL<312> A_IWL<311> A_IWL<310> A_IWL<309> A_IWL<308> A_IWL<307> A_IWL<306> A_IWL<305> A_IWL<304> A_IWL<303> A_IWL<302> A_IWL<301> A_IWL<300> A_IWL<299> A_IWL<298> A_IWL<297> A_IWL<296> A_IWL<295> A_IWL<294> A_IWL<293> A_IWL<292> A_IWL<291> A_IWL<290> A_IWL<289> A_IWL<288> A_IWL<287> A_IWL<286> A_IWL<285> A_IWL<284> A_IWL<283> A_IWL<282> A_IWL<281> A_IWL<280> A_IWL<279> A_IWL<278> A_IWL<277> A_IWL<276> A_IWL<275> A_IWL<274> A_IWL<273> A_IWL<272> A_IWL<271> A_IWL<270> A_IWL<269> A_IWL<268> A_IWL<267> A_IWL<266> A_IWL<265> A_IWL<264> A_IWL<263> A_IWL<262> A_IWL<261> A_IWL<260> A_IWL<259> A_IWL<258> A_IWL<257> A_IWL<256> A_IWL<255> A_IWL<254> A_IWL<253> A_IWL<252> A_IWL<251> A_IWL<250> A_IWL<249> A_IWL<248> A_IWL<247> A_IWL<246> A_IWL<245> A_IWL<244> A_IWL<243> A_IWL<242> A_IWL<241> A_IWL<240> A_IWL<239> A_IWL<238> A_IWL<237> A_IWL<236> A_IWL<235> A_IWL<234> A_IWL<233> A_IWL<232> A_IWL<231> A_IWL<230> A_IWL<229> A_IWL<228> A_IWL<227> A_IWL<226> A_IWL<225> A_IWL<224> A_IWL<223> A_IWL<222> A_IWL<221> A_IWL<220> A_IWL<219> A_IWL<218> A_IWL<217> A_IWL<216> A_IWL<215> A_IWL<214> A_IWL<213> A_IWL<212> A_IWL<211> A_IWL<210> A_IWL<209> A_IWL<208> A_IWL<207> A_IWL<206> A_IWL<205> A_IWL<204> A_IWL<203> A_IWL<202> A_IWL<201> A_IWL<200> A_IWL<199> A_IWL<198> A_IWL<197> A_IWL<196> A_IWL<195> A_IWL<194> A_IWL<193> A_IWL<192> A_IWL<191> A_IWL<190> A_IWL<189> A_IWL<188> A_IWL<187> A_IWL<186> A_IWL<185> A_IWL<184> A_IWL<183> A_IWL<182> A_IWL<181> A_IWL<180> A_IWL<179> A_IWL<178> A_IWL<177> A_IWL<176> A_IWL<175> A_IWL<174> A_IWL<173> A_IWL<172> A_IWL<171> A_IWL<170> A_IWL<169> A_IWL<168> A_IWL<167> A_IWL<166> A_IWL<165> A_IWL<164> A_IWL<163> A_IWL<162> A_IWL<161> A_IWL<160> A_IWL<159> A_IWL<158> A_IWL<157> A_IWL<156> A_IWL<155> A_IWL<154> A_IWL<153> A_IWL<152> A_IWL<151> A_IWL<150> A_IWL<149> A_IWL<148> A_IWL<147> A_IWL<146> A_IWL<145> A_IWL<144> A_IWL<143> A_IWL<142> A_IWL<141> A_IWL<140> A_IWL<139> A_IWL<138> A_IWL<137> A_IWL<136> A_IWL<135> A_IWL<134> A_IWL<133> A_IWL<132> A_IWL<131> A_IWL<130> A_IWL<129> A_IWL<128> A_IWL<127> A_IWL<126> A_IWL<125> A_IWL<124> A_IWL<123> A_IWL<122> A_IWL<121> A_IWL<120> A_IWL<119> A_IWL<118> A_IWL<117> A_IWL<116> A_IWL<115> A_IWL<114> A_IWL<113> A_IWL<112> A_IWL<111> A_IWL<110> A_IWL<109> A_IWL<108> A_IWL<107> A_IWL<106> A_IWL<105> A_IWL<104> A_IWL<103> A_IWL<102> A_IWL<101> A_IWL<100> A_IWL<99> A_IWL<98> A_IWL<97> A_IWL<96> A_IWL<95> A_IWL<94> A_IWL<93> A_IWL<92> A_IWL<91> A_IWL<90> A_IWL<89> A_IWL<88> A_IWL<87> A_IWL<86> A_IWL<85> A_IWL<84> A_IWL<83> A_IWL<82> A_IWL<81> A_IWL<80> A_IWL<79> A_IWL<78> A_IWL<77> A_IWL<76> A_IWL<75> A_IWL<74> A_IWL<73> A_IWL<72> A_IWL<71> A_IWL<70> A_IWL<69> A_IWL<68> A_IWL<67> A_IWL<66> A_IWL<65> A_IWL<64> A_IWL<63> A_IWL<62> A_IWL<61> A_IWL<60> A_IWL<59> A_IWL<58> A_IWL<57> A_IWL<56> A_IWL<55> A_IWL<54> A_IWL<53> A_IWL<52> A_IWL<51> A_IWL<50> A_IWL<49> A_IWL<48> A_IWL<47> A_IWL<46> A_IWL<45> A_IWL<44> A_IWL<43> A_IWL<42> A_IWL<41> A_IWL<40> A_IWL<39> A_IWL<38> A_IWL<37> A_IWL<36> A_IWL<35> A_IWL<34> A_IWL<33> A_IWL<32> A_IWL<31> A_IWL<30> A_IWL<29> A_IWL<28> A_IWL<27> A_IWL<26> A_IWL<25> A_IWL<24> A_IWL<23> A_IWL<22> A_IWL<21> A_IWL<20> A_IWL<19> A_IWL<18> A_IWL<17> A_IWL<16> A_IWL<15> A_IWL<14> A_IWL<13> A_IWL<12> A_IWL<11> A_IWL<10> A_IWL<9> A_IWL<8> A_IWL<7> A_IWL<6> A_IWL<5> A_IWL<4> A_IWL<3> A_IWL<2> A_IWL<1> A_IWL<0> VDD_CORE VSS / RM_IHPSG13_2048x64_c2_1P_COLUMN_pcell_0
.ENDS




.SUBCKT RM_IHPSG13_2048x64_c2_1P_DLY_pcell_2 A Z VDD VSS
	XIDL<3> D<7> Z VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<2> D<6> D<7> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<1> D<5> D<6> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDM<5> D<4> D<5> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<4> D<3> D<4> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<3> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<2> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
	XIDM<1> A D<1> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
.ENDS


.SUBCKT RM_IHPSG13_2048x64_c2_1P_DLY_pcell_3 A Z VDD VSS
	XIDL<7> D<7> Z VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<6> D<6> D<7> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<5> D<5> D<6> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<4> D<4> D<5> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<3> D<3> D<4> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<2> D<2> D<3> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDL<1> D<1> D<2> VDD VSS / RSC_IHPSG13_CDLYX1 
	XIDM A D<1> VDD VSS / RSC_IHPSG13_CDLYX1_DUMMY 
.ENDS



.SUBCKT RM_IHPSG13_1P_2048x64_c2_bm_bist A_ADDR<10> A_ADDR<9> A_ADDR<8> A_ADDR<7> A_ADDR<6> A_ADDR<5> A_ADDR<4> A_ADDR<3> A_ADDR<2> A_ADDR<1> A_ADDR<0> A_BIST_ADDR<10> A_BIST_ADDR<9> A_BIST_ADDR<8> A_BIST_ADDR<7> A_BIST_ADDR<6> A_BIST_ADDR<5> A_BIST_ADDR<4> A_BIST_ADDR<3> A_BIST_ADDR<2> A_BIST_ADDR<1> A_BIST_ADDR<0> A_BIST_BM<63> A_BIST_BM<62> A_BIST_BM<61> A_BIST_BM<60> A_BIST_BM<59> A_BIST_BM<58> A_BIST_BM<57> A_BIST_BM<56> A_BIST_BM<55> A_BIST_BM<54> A_BIST_BM<53> A_BIST_BM<52> A_BIST_BM<51> A_BIST_BM<50> A_BIST_BM<49> A_BIST_BM<48> A_BIST_BM<47> A_BIST_BM<46> A_BIST_BM<45> A_BIST_BM<44> A_BIST_BM<43> A_BIST_BM<42> A_BIST_BM<41> A_BIST_BM<40> A_BIST_BM<39> A_BIST_BM<38> A_BIST_BM<37> A_BIST_BM<36> A_BIST_BM<35> A_BIST_BM<34> A_BIST_BM<33> A_BIST_BM<32> A_BIST_BM<31> A_BIST_BM<30> A_BIST_BM<29> A_BIST_BM<28> A_BIST_BM<27> A_BIST_BM<26> A_BIST_BM<25> A_BIST_BM<24> A_BIST_BM<23> A_BIST_BM<22> A_BIST_BM<21> A_BIST_BM<20> A_BIST_BM<19> A_BIST_BM<18> A_BIST_BM<17> A_BIST_BM<16> A_BIST_BM<15> A_BIST_BM<14> A_BIST_BM<13> A_BIST_BM<12> A_BIST_BM<11> A_BIST_BM<10> A_BIST_BM<9> A_BIST_BM<8> A_BIST_BM<7> A_BIST_BM<6> A_BIST_BM<5> A_BIST_BM<4> A_BIST_BM<3> A_BIST_BM<2> A_BIST_BM<1> A_BIST_BM<0> A_BIST_CLK A_BIST_DIN<63> A_BIST_DIN<62> A_BIST_DIN<61> A_BIST_DIN<60> A_BIST_DIN<59> A_BIST_DIN<58> A_BIST_DIN<57> A_BIST_DIN<56> A_BIST_DIN<55> A_BIST_DIN<54> A_BIST_DIN<53> A_BIST_DIN<52> A_BIST_DIN<51> A_BIST_DIN<50> A_BIST_DIN<49> A_BIST_DIN<48> A_BIST_DIN<47> A_BIST_DIN<46> A_BIST_DIN<45> A_BIST_DIN<44> A_BIST_DIN<43> A_BIST_DIN<42> A_BIST_DIN<41> A_BIST_DIN<40> A_BIST_DIN<39> A_BIST_DIN<38> A_BIST_DIN<37> A_BIST_DIN<36> A_BIST_DIN<35> A_BIST_DIN<34> A_BIST_DIN<33> A_BIST_DIN<32> A_BIST_DIN<31> A_BIST_DIN<30> A_BIST_DIN<29> A_BIST_DIN<28> A_BIST_DIN<27> A_BIST_DIN<26> A_BIST_DIN<25> A_BIST_DIN<24> A_BIST_DIN<23> A_BIST_DIN<22> A_BIST_DIN<21> A_BIST_DIN<20> A_BIST_DIN<19> A_BIST_DIN<18> A_BIST_DIN<17> A_BIST_DIN<16> A_BIST_DIN<15> A_BIST_DIN<14> A_BIST_DIN<13> A_BIST_DIN<12> A_BIST_DIN<11> A_BIST_DIN<10> A_BIST_DIN<9> A_BIST_DIN<8> A_BIST_DIN<7> A_BIST_DIN<6> A_BIST_DIN<5> A_BIST_DIN<4> A_BIST_DIN<3> A_BIST_DIN<2> A_BIST_DIN<1> A_BIST_DIN<0> A_BIST_EN A_BIST_MEN A_BIST_REN A_BIST_WEN A_BM<63> A_BM<62> A_BM<61> A_BM<60> A_BM<59> A_BM<58> A_BM<57> A_BM<56> A_BM<55> A_BM<54> A_BM<53> A_BM<52> A_BM<51> A_BM<50> A_BM<49> A_BM<48> A_BM<47> A_BM<46> A_BM<45> A_BM<44> A_BM<43> A_BM<42> A_BM<41> A_BM<40> A_BM<39> A_BM<38> A_BM<37> A_BM<36> A_BM<35> A_BM<34> A_BM<33> A_BM<32> A_BM<31> A_BM<30> A_BM<29> A_BM<28> A_BM<27> A_BM<26> A_BM<25> A_BM<24> A_BM<23> A_BM<22> A_BM<21> A_BM<20> A_BM<19> A_BM<18> A_BM<17> A_BM<16> A_BM<15> A_BM<14> A_BM<13> A_BM<12> A_BM<11> A_BM<10> A_BM<9> A_BM<8> A_BM<7> A_BM<6> A_BM<5> A_BM<4> A_BM<3> A_BM<2> A_BM<1> A_BM<0> A_CLK A_DIN<63> A_DIN<62> A_DIN<61> A_DIN<60> A_DIN<59> A_DIN<58> A_DIN<57> A_DIN<56> A_DIN<55> A_DIN<54> A_DIN<53> A_DIN<52> A_DIN<51> A_DIN<50> A_DIN<49> A_DIN<48> A_DIN<47> A_DIN<46> A_DIN<45> A_DIN<44> A_DIN<43> A_DIN<42> A_DIN<41> A_DIN<40> A_DIN<39> A_DIN<38> A_DIN<37> A_DIN<36> A_DIN<35> A_DIN<34> A_DIN<33> A_DIN<32> A_DIN<31> A_DIN<30> A_DIN<29> A_DIN<28> A_DIN<27> A_DIN<26> A_DIN<25> A_DIN<24> A_DIN<23> A_DIN<22> A_DIN<21> A_DIN<20> A_DIN<19> A_DIN<18> A_DIN<17> A_DIN<16> A_DIN<15> A_DIN<14> A_DIN<13> A_DIN<12> A_DIN<11> A_DIN<10> A_DIN<9> A_DIN<8> A_DIN<7> A_DIN<6> A_DIN<5> A_DIN<4> A_DIN<3> A_DIN<2> A_DIN<1> A_DIN<0> A_DLY A_DOUT<63> A_DOUT<62> A_DOUT<61> A_DOUT<60> A_DOUT<59> A_DOUT<58> A_DOUT<57> A_DOUT<56> A_DOUT<55> A_DOUT<54> A_DOUT<53> A_DOUT<52> A_DOUT<51> A_DOUT<50> A_DOUT<49> A_DOUT<48> A_DOUT<47> A_DOUT<46> A_DOUT<45> A_DOUT<44> A_DOUT<43> A_DOUT<42> A_DOUT<41> A_DOUT<40> A_DOUT<39> A_DOUT<38> A_DOUT<37> A_DOUT<36> A_DOUT<35> A_DOUT<34> A_DOUT<33> A_DOUT<32> A_DOUT<31> A_DOUT<30> A_DOUT<29> A_DOUT<28> A_DOUT<27> A_DOUT<26> A_DOUT<25> A_DOUT<24> A_DOUT<23> A_DOUT<22> A_DOUT<21> A_DOUT<20> A_DOUT<19> A_DOUT<18> A_DOUT<17> A_DOUT<16> A_DOUT<15> A_DOUT<14> A_DOUT<13> A_DOUT<12> A_DOUT<11> A_DOUT<10> A_DOUT<9> A_DOUT<8> A_DOUT<7> A_DOUT<6> A_DOUT<5> A_DOUT<4> A_DOUT<3> A_DOUT<2> A_DOUT<1> A_DOUT<0> A_MEN A_REN A_WEN VDD! VDDARRAY! VSS!


XRAM<1> a_blc_r<127> a_blc_r<126> a_blc_r<125> a_blc_r<124> a_blc_r<123> a_blc_r<122> a_blc_r<121> a_blc_r<120> a_blc_r<119> a_blc_r<118> a_blc_r<117> a_blc_r<116> a_blc_r<115> a_blc_r<114> a_blc_r<113> a_blc_r<112> a_blc_r<111> a_blc_r<110> a_blc_r<109> a_blc_r<108> a_blc_r<107> a_blc_r<106> a_blc_r<105> a_blc_r<104> a_blc_r<103> a_blc_r<102> a_blc_r<101> a_blc_r<100> a_blc_r<99> a_blc_r<98> a_blc_r<97> a_blc_r<96> a_blc_r<95> a_blc_r<94> a_blc_r<93> a_blc_r<92> a_blc_r<91> a_blc_r<90> a_blc_r<89> a_blc_r<88> a_blc_r<87> a_blc_r<86> a_blc_r<85> a_blc_r<84> a_blc_r<83> a_blc_r<82> a_blc_r<81> a_blc_r<80> a_blc_r<79> a_blc_r<78> a_blc_r<77> a_blc_r<76> a_blc_r<75> a_blc_r<74> a_blc_r<73> a_blc_r<72> a_blc_r<71> a_blc_r<70> a_blc_r<69> a_blc_r<68> a_blc_r<67> a_blc_r<66> a_blc_r<65> a_blc_r<64> a_blc_r<63> a_blc_r<62> a_blc_r<61> a_blc_r<60> a_blc_r<59> a_blc_r<58> a_blc_r<57> a_blc_r<56> a_blc_r<55> a_blc_r<54> a_blc_r<53> a_blc_r<52> a_blc_r<51> a_blc_r<50> a_blc_r<49> a_blc_r<48> a_blc_r<47> a_blc_r<46> a_blc_r<45> a_blc_r<44> a_blc_r<43> a_blc_r<42> a_blc_r<41> a_blc_r<40> a_blc_r<39> a_blc_r<38> a_blc_r<37> a_blc_r<36> a_blc_r<35> a_blc_r<34> a_blc_r<33> a_blc_r<32> a_blc_r<31> a_blc_r<30> a_blc_r<29> a_blc_r<28> a_blc_r<27> a_blc_r<26> a_blc_r<25> a_blc_r<24> a_blc_r<23> a_blc_r<22> a_blc_r<21> a_blc_r<20> a_blc_r<19> a_blc_r<18> a_blc_r<17> a_blc_r<16> a_blc_r<15> a_blc_r<14> a_blc_r<13> a_blc_r<12> a_blc_r<11> a_blc_r<10> a_blc_r<9> a_blc_r<8> a_blc_r<7> a_blc_r<6> a_blc_r<5> a_blc_r<4> a_blc_r<3> a_blc_r<2> a_blc_r<1> a_blc_r<0> a_blt_r<127> a_blt_r<126> a_blt_r<125> a_blt_r<124> a_blt_r<123> a_blt_r<122> a_blt_r<121> a_blt_r<120> a_blt_r<119> a_blt_r<118> a_blt_r<117> a_blt_r<116> a_blt_r<115> a_blt_r<114> a_blt_r<113> a_blt_r<112> a_blt_r<111> a_blt_r<110> a_blt_r<109> a_blt_r<108> a_blt_r<107> a_blt_r<106> a_blt_r<105> a_blt_r<104> a_blt_r<103> a_blt_r<102> a_blt_r<101> a_blt_r<100> a_blt_r<99> a_blt_r<98> a_blt_r<97> a_blt_r<96> a_blt_r<95> a_blt_r<94> a_blt_r<93> a_blt_r<92> a_blt_r<91> a_blt_r<90> a_blt_r<89> a_blt_r<88> a_blt_r<87> a_blt_r<86> a_blt_r<85> a_blt_r<84> a_blt_r<83> a_blt_r<82> a_blt_r<81> a_blt_r<80> a_blt_r<79> a_blt_r<78> a_blt_r<77> a_blt_r<76> a_blt_r<75> a_blt_r<74> a_blt_r<73> a_blt_r<72> a_blt_r<71> a_blt_r<70> a_blt_r<69> a_blt_r<68> a_blt_r<67> a_blt_r<66> a_blt_r<65> a_blt_r<64> a_blt_r<63> a_blt_r<62> a_blt_r<61> a_blt_r<60> a_blt_r<59> a_blt_r<58> a_blt_r<57> a_blt_r<56> a_blt_r<55> a_blt_r<54> a_blt_r<53> a_blt_r<52> a_blt_r<51> a_blt_r<50> a_blt_r<49> a_blt_r<48> a_blt_r<47> a_blt_r<46> a_blt_r<45> a_blt_r<44> a_blt_r<43> a_blt_r<42> a_blt_r<41> a_blt_r<40> a_blt_r<39> a_blt_r<38> a_blt_r<37> a_blt_r<36> a_blt_r<35> a_blt_r<34> a_blt_r<33> a_blt_r<32> a_blt_r<31> a_blt_r<30> a_blt_r<29> a_blt_r<28> a_blt_r<27> a_blt_r<26> a_blt_r<25> a_blt_r<24> a_blt_r<23> a_blt_r<22> a_blt_r<21> a_blt_r<20> a_blt_r<19> a_blt_r<18> a_blt_r<17> a_blt_r<16> a_blt_r<15> a_blt_r<14> a_blt_r<13> a_blt_r<12> a_blt_r<11> a_blt_r<10> a_blt_r<9> a_blt_r<8> a_blt_r<7> a_blt_r<6> a_blt_r<5> a_blt_r<4> a_blt_r<3> a_blt_r<2> a_blt_r<1> a_blt_r<0> a_wl_r<511> a_wl_r<510> a_wl_r<509> a_wl_r<508> a_wl_r<507> a_wl_r<506> a_wl_r<505> a_wl_r<504> a_wl_r<503> a_wl_r<502> a_wl_r<501> a_wl_r<500> a_wl_r<499> a_wl_r<498> a_wl_r<497> a_wl_r<496> a_wl_r<495> a_wl_r<494> a_wl_r<493> a_wl_r<492> a_wl_r<491> a_wl_r<490> a_wl_r<489> a_wl_r<488> a_wl_r<487> a_wl_r<486> a_wl_r<485> a_wl_r<484> a_wl_r<483> a_wl_r<482> a_wl_r<481> a_wl_r<480> a_wl_r<479> a_wl_r<478> a_wl_r<477> a_wl_r<476> a_wl_r<475> a_wl_r<474> a_wl_r<473> a_wl_r<472> a_wl_r<471> a_wl_r<470> a_wl_r<469> a_wl_r<468> a_wl_r<467> a_wl_r<466> a_wl_r<465> a_wl_r<464> a_wl_r<463> a_wl_r<462> a_wl_r<461> a_wl_r<460> a_wl_r<459> a_wl_r<458> a_wl_r<457> a_wl_r<456> a_wl_r<455> a_wl_r<454> a_wl_r<453> a_wl_r<452> a_wl_r<451> a_wl_r<450> a_wl_r<449> a_wl_r<448> a_wl_r<447> a_wl_r<446> a_wl_r<445> a_wl_r<444> a_wl_r<443> a_wl_r<442> a_wl_r<441> a_wl_r<440> a_wl_r<439> a_wl_r<438> a_wl_r<437> a_wl_r<436> a_wl_r<435> a_wl_r<434> a_wl_r<433> a_wl_r<432> a_wl_r<431> a_wl_r<430> a_wl_r<429> a_wl_r<428> a_wl_r<427> a_wl_r<426> a_wl_r<425> a_wl_r<424> a_wl_r<423> a_wl_r<422> a_wl_r<421> a_wl_r<420> a_wl_r<419> a_wl_r<418> a_wl_r<417> a_wl_r<416> a_wl_r<415> a_wl_r<414> a_wl_r<413> a_wl_r<412> a_wl_r<411> a_wl_r<410> a_wl_r<409> a_wl_r<408> a_wl_r<407> a_wl_r<406> a_wl_r<405> a_wl_r<404> a_wl_r<403> a_wl_r<402> a_wl_r<401> a_wl_r<400> a_wl_r<399> a_wl_r<398> a_wl_r<397> a_wl_r<396> a_wl_r<395> a_wl_r<394> a_wl_r<393> a_wl_r<392> a_wl_r<391> a_wl_r<390> a_wl_r<389> a_wl_r<388> a_wl_r<387> a_wl_r<386> a_wl_r<385> a_wl_r<384> a_wl_r<383> a_wl_r<382> a_wl_r<381> a_wl_r<380> a_wl_r<379> a_wl_r<378> a_wl_r<377> a_wl_r<376> a_wl_r<375> a_wl_r<374> a_wl_r<373> a_wl_r<372> a_wl_r<371> a_wl_r<370> a_wl_r<369> a_wl_r<368> a_wl_r<367> a_wl_r<366> a_wl_r<365> a_wl_r<364> a_wl_r<363> a_wl_r<362> a_wl_r<361> a_wl_r<360> a_wl_r<359> a_wl_r<358> a_wl_r<357> a_wl_r<356> a_wl_r<355> a_wl_r<354> a_wl_r<353> a_wl_r<352> a_wl_r<351> a_wl_r<350> a_wl_r<349> a_wl_r<348> a_wl_r<347> a_wl_r<346> a_wl_r<345> a_wl_r<344> a_wl_r<343> a_wl_r<342> a_wl_r<341> a_wl_r<340> a_wl_r<339> a_wl_r<338> a_wl_r<337> a_wl_r<336> a_wl_r<335> a_wl_r<334> a_wl_r<333> a_wl_r<332> a_wl_r<331> a_wl_r<330> a_wl_r<329> a_wl_r<328> a_wl_r<327> a_wl_r<326> a_wl_r<325> a_wl_r<324> a_wl_r<323> a_wl_r<322> a_wl_r<321> a_wl_r<320> a_wl_r<319> a_wl_r<318> a_wl_r<317> a_wl_r<316> a_wl_r<315> a_wl_r<314> a_wl_r<313> a_wl_r<312> a_wl_r<311> a_wl_r<310> a_wl_r<309> a_wl_r<308> a_wl_r<307> a_wl_r<306> a_wl_r<305> a_wl_r<304> a_wl_r<303> a_wl_r<302> a_wl_r<301> a_wl_r<300> a_wl_r<299> a_wl_r<298> a_wl_r<297> a_wl_r<296> a_wl_r<295> a_wl_r<294> a_wl_r<293> a_wl_r<292> a_wl_r<291> a_wl_r<290> a_wl_r<289> a_wl_r<288> a_wl_r<287> a_wl_r<286> a_wl_r<285> a_wl_r<284> a_wl_r<283> a_wl_r<282> a_wl_r<281> a_wl_r<280> a_wl_r<279> a_wl_r<278> a_wl_r<277> a_wl_r<276> a_wl_r<275> a_wl_r<274> a_wl_r<273> a_wl_r<272> a_wl_r<271> a_wl_r<270> a_wl_r<269> a_wl_r<268> a_wl_r<267> a_wl_r<266> a_wl_r<265> a_wl_r<264> a_wl_r<263> a_wl_r<262> a_wl_r<261> a_wl_r<260> a_wl_r<259> a_wl_r<258> a_wl_r<257> a_wl_r<256> a_wl_r<255> a_wl_r<254> a_wl_r<253> a_wl_r<252> a_wl_r<251> a_wl_r<250> a_wl_r<249> a_wl_r<248> a_wl_r<247> a_wl_r<246> a_wl_r<245> a_wl_r<244> a_wl_r<243> a_wl_r<242> a_wl_r<241> a_wl_r<240> a_wl_r<239> a_wl_r<238> a_wl_r<237> a_wl_r<236> a_wl_r<235> a_wl_r<234> a_wl_r<233> a_wl_r<232> a_wl_r<231> a_wl_r<230> a_wl_r<229> a_wl_r<228> a_wl_r<227> a_wl_r<226> a_wl_r<225> a_wl_r<224> a_wl_r<223> a_wl_r<222> a_wl_r<221> a_wl_r<220> a_wl_r<219> a_wl_r<218> a_wl_r<217> a_wl_r<216> a_wl_r<215> a_wl_r<214> a_wl_r<213> a_wl_r<212> a_wl_r<211> a_wl_r<210> a_wl_r<209> a_wl_r<208> a_wl_r<207> a_wl_r<206> a_wl_r<205> a_wl_r<204> a_wl_r<203> a_wl_r<202> a_wl_r<201> a_wl_r<200> a_wl_r<199> a_wl_r<198> a_wl_r<197> a_wl_r<196> a_wl_r<195> a_wl_r<194> a_wl_r<193> a_wl_r<192> a_wl_r<191> a_wl_r<190> a_wl_r<189> a_wl_r<188> a_wl_r<187> a_wl_r<186> a_wl_r<185> a_wl_r<184> a_wl_r<183> a_wl_r<182> a_wl_r<181> a_wl_r<180> a_wl_r<179> a_wl_r<178> a_wl_r<177> a_wl_r<176> a_wl_r<175> a_wl_r<174> a_wl_r<173> a_wl_r<172> a_wl_r<171> a_wl_r<170> a_wl_r<169> a_wl_r<168> a_wl_r<167> a_wl_r<166> a_wl_r<165> a_wl_r<164> a_wl_r<163> a_wl_r<162> a_wl_r<161> a_wl_r<160> a_wl_r<159> a_wl_r<158> a_wl_r<157> a_wl_r<156> a_wl_r<155> a_wl_r<154> a_wl_r<153> a_wl_r<152> a_wl_r<151> a_wl_r<150> a_wl_r<149> a_wl_r<148> a_wl_r<147> a_wl_r<146> a_wl_r<145> a_wl_r<144> a_wl_r<143> a_wl_r<142> a_wl_r<141> a_wl_r<140> a_wl_r<139> a_wl_r<138> a_wl_r<137> a_wl_r<136> a_wl_r<135> a_wl_r<134> a_wl_r<133> a_wl_r<132> a_wl_r<131> a_wl_r<130> a_wl_r<129> a_wl_r<128> a_wl_r<127> a_wl_r<126> a_wl_r<125> a_wl_r<124> a_wl_r<123> a_wl_r<122> a_wl_r<121> a_wl_r<120> a_wl_r<119> a_wl_r<118> a_wl_r<117> a_wl_r<116> a_wl_r<115> a_wl_r<114> a_wl_r<113> a_wl_r<112> a_wl_r<111> a_wl_r<110> a_wl_r<109> a_wl_r<108> a_wl_r<107> a_wl_r<106> a_wl_r<105> a_wl_r<104> a_wl_r<103> a_wl_r<102> a_wl_r<101> a_wl_r<100> a_wl_r<99> a_wl_r<98> a_wl_r<97> a_wl_r<96> a_wl_r<95> a_wl_r<94> a_wl_r<93> a_wl_r<92> a_wl_r<91> a_wl_r<90> a_wl_r<89> a_wl_r<88> a_wl_r<87> a_wl_r<86> a_wl_r<85> a_wl_r<84> a_wl_r<83> a_wl_r<82> a_wl_r<81> a_wl_r<80> a_wl_r<79> a_wl_r<78> a_wl_r<77> a_wl_r<76> a_wl_r<75> a_wl_r<74> a_wl_r<73> a_wl_r<72> a_wl_r<71> a_wl_r<70> a_wl_r<69> a_wl_r<68> a_wl_r<67> a_wl_r<66> a_wl_r<65> a_wl_r<64> a_wl_r<63> a_wl_r<62> a_wl_r<61> a_wl_r<60> a_wl_r<59> a_wl_r<58> a_wl_r<57> a_wl_r<56> a_wl_r<55> a_wl_r<54> a_wl_r<53> a_wl_r<52> a_wl_r<51> a_wl_r<50> a_wl_r<49> a_wl_r<48> a_wl_r<47> a_wl_r<46> a_wl_r<45> a_wl_r<44> a_wl_r<43> a_wl_r<42> a_wl_r<41> a_wl_r<40> a_wl_r<39> a_wl_r<38> a_wl_r<37> a_wl_r<36> a_wl_r<35> a_wl_r<34> a_wl_r<33> a_wl_r<32> a_wl_r<31> a_wl_r<30> a_wl_r<29> a_wl_r<28> a_wl_r<27> a_wl_r<26> a_wl_r<25> a_wl_r<24> a_wl_r<23> a_wl_r<22> a_wl_r<21> a_wl_r<20> a_wl_r<19> a_wl_r<18> a_wl_r<17> a_wl_r<16> a_wl_r<15> a_wl_r<14> a_wl_r<13> a_wl_r<12> a_wl_r<11> a_wl_r<10> a_wl_r<9> a_wl_r<8> a_wl_r<7> a_wl_r<6> a_wl_r<5> a_wl_r<4> a_wl_r<3> a_wl_r<2> a_wl_r<1> a_wl_r<0> VDDARRAY! VSS! / RM_IHPSG13_2048x64_c2_1P_MATRIX_pcell_1
XRAM<0> a_blc_l<127> a_blc_l<126> a_blc_l<125> a_blc_l<124> a_blc_l<123> a_blc_l<122> a_blc_l<121> a_blc_l<120> a_blc_l<119> a_blc_l<118> a_blc_l<117> a_blc_l<116> a_blc_l<115> a_blc_l<114> a_blc_l<113> a_blc_l<112> a_blc_l<111> a_blc_l<110> a_blc_l<109> a_blc_l<108> a_blc_l<107> a_blc_l<106> a_blc_l<105> a_blc_l<104> a_blc_l<103> a_blc_l<102> a_blc_l<101> a_blc_l<100> a_blc_l<99> a_blc_l<98> a_blc_l<97> a_blc_l<96> a_blc_l<95> a_blc_l<94> a_blc_l<93> a_blc_l<92> a_blc_l<91> a_blc_l<90> a_blc_l<89> a_blc_l<88> a_blc_l<87> a_blc_l<86> a_blc_l<85> a_blc_l<84> a_blc_l<83> a_blc_l<82> a_blc_l<81> a_blc_l<80> a_blc_l<79> a_blc_l<78> a_blc_l<77> a_blc_l<76> a_blc_l<75> a_blc_l<74> a_blc_l<73> a_blc_l<72> a_blc_l<71> a_blc_l<70> a_blc_l<69> a_blc_l<68> a_blc_l<67> a_blc_l<66> a_blc_l<65> a_blc_l<64> a_blc_l<63> a_blc_l<62> a_blc_l<61> a_blc_l<60> a_blc_l<59> a_blc_l<58> a_blc_l<57> a_blc_l<56> a_blc_l<55> a_blc_l<54> a_blc_l<53> a_blc_l<52> a_blc_l<51> a_blc_l<50> a_blc_l<49> a_blc_l<48> a_blc_l<47> a_blc_l<46> a_blc_l<45> a_blc_l<44> a_blc_l<43> a_blc_l<42> a_blc_l<41> a_blc_l<40> a_blc_l<39> a_blc_l<38> a_blc_l<37> a_blc_l<36> a_blc_l<35> a_blc_l<34> a_blc_l<33> a_blc_l<32> a_blc_l<31> a_blc_l<30> a_blc_l<29> a_blc_l<28> a_blc_l<27> a_blc_l<26> a_blc_l<25> a_blc_l<24> a_blc_l<23> a_blc_l<22> a_blc_l<21> a_blc_l<20> a_blc_l<19> a_blc_l<18> a_blc_l<17> a_blc_l<16> a_blc_l<15> a_blc_l<14> a_blc_l<13> a_blc_l<12> a_blc_l<11> a_blc_l<10> a_blc_l<9> a_blc_l<8> a_blc_l<7> a_blc_l<6> a_blc_l<5> a_blc_l<4> a_blc_l<3> a_blc_l<2> a_blc_l<1> a_blc_l<0> a_blt_l<127> a_blt_l<126> a_blt_l<125> a_blt_l<124> a_blt_l<123> a_blt_l<122> a_blt_l<121> a_blt_l<120> a_blt_l<119> a_blt_l<118> a_blt_l<117> a_blt_l<116> a_blt_l<115> a_blt_l<114> a_blt_l<113> a_blt_l<112> a_blt_l<111> a_blt_l<110> a_blt_l<109> a_blt_l<108> a_blt_l<107> a_blt_l<106> a_blt_l<105> a_blt_l<104> a_blt_l<103> a_blt_l<102> a_blt_l<101> a_blt_l<100> a_blt_l<99> a_blt_l<98> a_blt_l<97> a_blt_l<96> a_blt_l<95> a_blt_l<94> a_blt_l<93> a_blt_l<92> a_blt_l<91> a_blt_l<90> a_blt_l<89> a_blt_l<88> a_blt_l<87> a_blt_l<86> a_blt_l<85> a_blt_l<84> a_blt_l<83> a_blt_l<82> a_blt_l<81> a_blt_l<80> a_blt_l<79> a_blt_l<78> a_blt_l<77> a_blt_l<76> a_blt_l<75> a_blt_l<74> a_blt_l<73> a_blt_l<72> a_blt_l<71> a_blt_l<70> a_blt_l<69> a_blt_l<68> a_blt_l<67> a_blt_l<66> a_blt_l<65> a_blt_l<64> a_blt_l<63> a_blt_l<62> a_blt_l<61> a_blt_l<60> a_blt_l<59> a_blt_l<58> a_blt_l<57> a_blt_l<56> a_blt_l<55> a_blt_l<54> a_blt_l<53> a_blt_l<52> a_blt_l<51> a_blt_l<50> a_blt_l<49> a_blt_l<48> a_blt_l<47> a_blt_l<46> a_blt_l<45> a_blt_l<44> a_blt_l<43> a_blt_l<42> a_blt_l<41> a_blt_l<40> a_blt_l<39> a_blt_l<38> a_blt_l<37> a_blt_l<36> a_blt_l<35> a_blt_l<34> a_blt_l<33> a_blt_l<32> a_blt_l<31> a_blt_l<30> a_blt_l<29> a_blt_l<28> a_blt_l<27> a_blt_l<26> a_blt_l<25> a_blt_l<24> a_blt_l<23> a_blt_l<22> a_blt_l<21> a_blt_l<20> a_blt_l<19> a_blt_l<18> a_blt_l<17> a_blt_l<16> a_blt_l<15> a_blt_l<14> a_blt_l<13> a_blt_l<12> a_blt_l<11> a_blt_l<10> a_blt_l<9> a_blt_l<8> a_blt_l<7> a_blt_l<6> a_blt_l<5> a_blt_l<4> a_blt_l<3> a_blt_l<2> a_blt_l<1> a_blt_l<0> a_wl_l<511> a_wl_l<510> a_wl_l<509> a_wl_l<508> a_wl_l<507> a_wl_l<506> a_wl_l<505> a_wl_l<504> a_wl_l<503> a_wl_l<502> a_wl_l<501> a_wl_l<500> a_wl_l<499> a_wl_l<498> a_wl_l<497> a_wl_l<496> a_wl_l<495> a_wl_l<494> a_wl_l<493> a_wl_l<492> a_wl_l<491> a_wl_l<490> a_wl_l<489> a_wl_l<488> a_wl_l<487> a_wl_l<486> a_wl_l<485> a_wl_l<484> a_wl_l<483> a_wl_l<482> a_wl_l<481> a_wl_l<480> a_wl_l<479> a_wl_l<478> a_wl_l<477> a_wl_l<476> a_wl_l<475> a_wl_l<474> a_wl_l<473> a_wl_l<472> a_wl_l<471> a_wl_l<470> a_wl_l<469> a_wl_l<468> a_wl_l<467> a_wl_l<466> a_wl_l<465> a_wl_l<464> a_wl_l<463> a_wl_l<462> a_wl_l<461> a_wl_l<460> a_wl_l<459> a_wl_l<458> a_wl_l<457> a_wl_l<456> a_wl_l<455> a_wl_l<454> a_wl_l<453> a_wl_l<452> a_wl_l<451> a_wl_l<450> a_wl_l<449> a_wl_l<448> a_wl_l<447> a_wl_l<446> a_wl_l<445> a_wl_l<444> a_wl_l<443> a_wl_l<442> a_wl_l<441> a_wl_l<440> a_wl_l<439> a_wl_l<438> a_wl_l<437> a_wl_l<436> a_wl_l<435> a_wl_l<434> a_wl_l<433> a_wl_l<432> a_wl_l<431> a_wl_l<430> a_wl_l<429> a_wl_l<428> a_wl_l<427> a_wl_l<426> a_wl_l<425> a_wl_l<424> a_wl_l<423> a_wl_l<422> a_wl_l<421> a_wl_l<420> a_wl_l<419> a_wl_l<418> a_wl_l<417> a_wl_l<416> a_wl_l<415> a_wl_l<414> a_wl_l<413> a_wl_l<412> a_wl_l<411> a_wl_l<410> a_wl_l<409> a_wl_l<408> a_wl_l<407> a_wl_l<406> a_wl_l<405> a_wl_l<404> a_wl_l<403> a_wl_l<402> a_wl_l<401> a_wl_l<400> a_wl_l<399> a_wl_l<398> a_wl_l<397> a_wl_l<396> a_wl_l<395> a_wl_l<394> a_wl_l<393> a_wl_l<392> a_wl_l<391> a_wl_l<390> a_wl_l<389> a_wl_l<388> a_wl_l<387> a_wl_l<386> a_wl_l<385> a_wl_l<384> a_wl_l<383> a_wl_l<382> a_wl_l<381> a_wl_l<380> a_wl_l<379> a_wl_l<378> a_wl_l<377> a_wl_l<376> a_wl_l<375> a_wl_l<374> a_wl_l<373> a_wl_l<372> a_wl_l<371> a_wl_l<370> a_wl_l<369> a_wl_l<368> a_wl_l<367> a_wl_l<366> a_wl_l<365> a_wl_l<364> a_wl_l<363> a_wl_l<362> a_wl_l<361> a_wl_l<360> a_wl_l<359> a_wl_l<358> a_wl_l<357> a_wl_l<356> a_wl_l<355> a_wl_l<354> a_wl_l<353> a_wl_l<352> a_wl_l<351> a_wl_l<350> a_wl_l<349> a_wl_l<348> a_wl_l<347> a_wl_l<346> a_wl_l<345> a_wl_l<344> a_wl_l<343> a_wl_l<342> a_wl_l<341> a_wl_l<340> a_wl_l<339> a_wl_l<338> a_wl_l<337> a_wl_l<336> a_wl_l<335> a_wl_l<334> a_wl_l<333> a_wl_l<332> a_wl_l<331> a_wl_l<330> a_wl_l<329> a_wl_l<328> a_wl_l<327> a_wl_l<326> a_wl_l<325> a_wl_l<324> a_wl_l<323> a_wl_l<322> a_wl_l<321> a_wl_l<320> a_wl_l<319> a_wl_l<318> a_wl_l<317> a_wl_l<316> a_wl_l<315> a_wl_l<314> a_wl_l<313> a_wl_l<312> a_wl_l<311> a_wl_l<310> a_wl_l<309> a_wl_l<308> a_wl_l<307> a_wl_l<306> a_wl_l<305> a_wl_l<304> a_wl_l<303> a_wl_l<302> a_wl_l<301> a_wl_l<300> a_wl_l<299> a_wl_l<298> a_wl_l<297> a_wl_l<296> a_wl_l<295> a_wl_l<294> a_wl_l<293> a_wl_l<292> a_wl_l<291> a_wl_l<290> a_wl_l<289> a_wl_l<288> a_wl_l<287> a_wl_l<286> a_wl_l<285> a_wl_l<284> a_wl_l<283> a_wl_l<282> a_wl_l<281> a_wl_l<280> a_wl_l<279> a_wl_l<278> a_wl_l<277> a_wl_l<276> a_wl_l<275> a_wl_l<274> a_wl_l<273> a_wl_l<272> a_wl_l<271> a_wl_l<270> a_wl_l<269> a_wl_l<268> a_wl_l<267> a_wl_l<266> a_wl_l<265> a_wl_l<264> a_wl_l<263> a_wl_l<262> a_wl_l<261> a_wl_l<260> a_wl_l<259> a_wl_l<258> a_wl_l<257> a_wl_l<256> a_wl_l<255> a_wl_l<254> a_wl_l<253> a_wl_l<252> a_wl_l<251> a_wl_l<250> a_wl_l<249> a_wl_l<248> a_wl_l<247> a_wl_l<246> a_wl_l<245> a_wl_l<244> a_wl_l<243> a_wl_l<242> a_wl_l<241> a_wl_l<240> a_wl_l<239> a_wl_l<238> a_wl_l<237> a_wl_l<236> a_wl_l<235> a_wl_l<234> a_wl_l<233> a_wl_l<232> a_wl_l<231> a_wl_l<230> a_wl_l<229> a_wl_l<228> a_wl_l<227> a_wl_l<226> a_wl_l<225> a_wl_l<224> a_wl_l<223> a_wl_l<222> a_wl_l<221> a_wl_l<220> a_wl_l<219> a_wl_l<218> a_wl_l<217> a_wl_l<216> a_wl_l<215> a_wl_l<214> a_wl_l<213> a_wl_l<212> a_wl_l<211> a_wl_l<210> a_wl_l<209> a_wl_l<208> a_wl_l<207> a_wl_l<206> a_wl_l<205> a_wl_l<204> a_wl_l<203> a_wl_l<202> a_wl_l<201> a_wl_l<200> a_wl_l<199> a_wl_l<198> a_wl_l<197> a_wl_l<196> a_wl_l<195> a_wl_l<194> a_wl_l<193> a_wl_l<192> a_wl_l<191> a_wl_l<190> a_wl_l<189> a_wl_l<188> a_wl_l<187> a_wl_l<186> a_wl_l<185> a_wl_l<184> a_wl_l<183> a_wl_l<182> a_wl_l<181> a_wl_l<180> a_wl_l<179> a_wl_l<178> a_wl_l<177> a_wl_l<176> a_wl_l<175> a_wl_l<174> a_wl_l<173> a_wl_l<172> a_wl_l<171> a_wl_l<170> a_wl_l<169> a_wl_l<168> a_wl_l<167> a_wl_l<166> a_wl_l<165> a_wl_l<164> a_wl_l<163> a_wl_l<162> a_wl_l<161> a_wl_l<160> a_wl_l<159> a_wl_l<158> a_wl_l<157> a_wl_l<156> a_wl_l<155> a_wl_l<154> a_wl_l<153> a_wl_l<152> a_wl_l<151> a_wl_l<150> a_wl_l<149> a_wl_l<148> a_wl_l<147> a_wl_l<146> a_wl_l<145> a_wl_l<144> a_wl_l<143> a_wl_l<142> a_wl_l<141> a_wl_l<140> a_wl_l<139> a_wl_l<138> a_wl_l<137> a_wl_l<136> a_wl_l<135> a_wl_l<134> a_wl_l<133> a_wl_l<132> a_wl_l<131> a_wl_l<130> a_wl_l<129> a_wl_l<128> a_wl_l<127> a_wl_l<126> a_wl_l<125> a_wl_l<124> a_wl_l<123> a_wl_l<122> a_wl_l<121> a_wl_l<120> a_wl_l<119> a_wl_l<118> a_wl_l<117> a_wl_l<116> a_wl_l<115> a_wl_l<114> a_wl_l<113> a_wl_l<112> a_wl_l<111> a_wl_l<110> a_wl_l<109> a_wl_l<108> a_wl_l<107> a_wl_l<106> a_wl_l<105> a_wl_l<104> a_wl_l<103> a_wl_l<102> a_wl_l<101> a_wl_l<100> a_wl_l<99> a_wl_l<98> a_wl_l<97> a_wl_l<96> a_wl_l<95> a_wl_l<94> a_wl_l<93> a_wl_l<92> a_wl_l<91> a_wl_l<90> a_wl_l<89> a_wl_l<88> a_wl_l<87> a_wl_l<86> a_wl_l<85> a_wl_l<84> a_wl_l<83> a_wl_l<82> a_wl_l<81> a_wl_l<80> a_wl_l<79> a_wl_l<78> a_wl_l<77> a_wl_l<76> a_wl_l<75> a_wl_l<74> a_wl_l<73> a_wl_l<72> a_wl_l<71> a_wl_l<70> a_wl_l<69> a_wl_l<68> a_wl_l<67> a_wl_l<66> a_wl_l<65> a_wl_l<64> a_wl_l<63> a_wl_l<62> a_wl_l<61> a_wl_l<60> a_wl_l<59> a_wl_l<58> a_wl_l<57> a_wl_l<56> a_wl_l<55> a_wl_l<54> a_wl_l<53> a_wl_l<52> a_wl_l<51> a_wl_l<50> a_wl_l<49> a_wl_l<48> a_wl_l<47> a_wl_l<46> a_wl_l<45> a_wl_l<44> a_wl_l<43> a_wl_l<42> a_wl_l<41> a_wl_l<40> a_wl_l<39> a_wl_l<38> a_wl_l<37> a_wl_l<36> a_wl_l<35> a_wl_l<34> a_wl_l<33> a_wl_l<32> a_wl_l<31> a_wl_l<30> a_wl_l<29> a_wl_l<28> a_wl_l<27> a_wl_l<26> a_wl_l<25> a_wl_l<24> a_wl_l<23> a_wl_l<22> a_wl_l<21> a_wl_l<20> a_wl_l<19> a_wl_l<18> a_wl_l<17> a_wl_l<16> a_wl_l<15> a_wl_l<14> a_wl_l<13> a_wl_l<12> a_wl_l<11> a_wl_l<10> a_wl_l<9> a_wl_l<8> a_wl_l<7> a_wl_l<6> a_wl_l<5> a_wl_l<4> a_wl_l<3> a_wl_l<2> a_wl_l<1> a_wl_l<0> VDDARRAY! VSS! / RM_IHPSG13_2048x64_c2_1P_MATRIX_pcell_1


XA_COLDRV<1> a_addr_col<1> a_addr_col<0> a_addr_col_r<1> a_addr_col_r<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> a_addr_dec_r<7> a_addr_dec_r<6> a_addr_dec_r<5> a_addr_dec_r<4> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> a_dclk a_dclk_p_r<0> a_rclk a_rclk_p_r<0> a_wclk a_wclk_p_r<0> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13X8
XA_COLDRV<0> a_addr_col<1> a_addr_col<0> a_addr_col_l<1> a_addr_col_l<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> a_addr_dec_l<7> a_addr_dec_l<6> a_addr_dec_l<5> a_addr_dec_l<4> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> a_dclk a_dclk_p_l<0> a_rclk a_rclk_p_l<0> a_wclk a_wclk_p_l<0> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13X8


XA_WLDRV<63> a_wi<511> a_wi<510> a_wi<509> a_wi<508> a_wi<507> a_wi<506> a_wi<505> a_wi<504> a_wi<503> a_wi<502> a_wi<501> a_wi<500> a_wi<499> a_wi<498> a_wi<497> a_wi<496> a_wl_r<511> a_wl_r<510> a_wl_r<509> a_wl_r<508> a_wl_r<507> a_wl_r<506> a_wl_r<505> a_wl_r<504> a_wl_r<503> a_wl_r<502> a_wl_r<501> a_wl_r<500> a_wl_r<499> a_wl_r<498> a_wl_r<497> a_wl_r<496>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<62> a_wi<495> a_wi<494> a_wi<493> a_wi<492> a_wi<491> a_wi<490> a_wi<489> a_wi<488> a_wi<487> a_wi<486> a_wi<485> a_wi<484> a_wi<483> a_wi<482> a_wi<481> a_wi<480> a_wl_r<495> a_wl_r<494> a_wl_r<493> a_wl_r<492> a_wl_r<491> a_wl_r<490> a_wl_r<489> a_wl_r<488> a_wl_r<487> a_wl_r<486> a_wl_r<485> a_wl_r<484> a_wl_r<483> a_wl_r<482> a_wl_r<481> a_wl_r<480>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<61> a_wi<479> a_wi<478> a_wi<477> a_wi<476> a_wi<475> a_wi<474> a_wi<473> a_wi<472> a_wi<471> a_wi<470> a_wi<469> a_wi<468> a_wi<467> a_wi<466> a_wi<465> a_wi<464> a_wl_r<479> a_wl_r<478> a_wl_r<477> a_wl_r<476> a_wl_r<475> a_wl_r<474> a_wl_r<473> a_wl_r<472> a_wl_r<471> a_wl_r<470> a_wl_r<469> a_wl_r<468> a_wl_r<467> a_wl_r<466> a_wl_r<465> a_wl_r<464>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<60> a_wi<463> a_wi<462> a_wi<461> a_wi<460> a_wi<459> a_wi<458> a_wi<457> a_wi<456> a_wi<455> a_wi<454> a_wi<453> a_wi<452> a_wi<451> a_wi<450> a_wi<449> a_wi<448> a_wl_r<463> a_wl_r<462> a_wl_r<461> a_wl_r<460> a_wl_r<459> a_wl_r<458> a_wl_r<457> a_wl_r<456> a_wl_r<455> a_wl_r<454> a_wl_r<453> a_wl_r<452> a_wl_r<451> a_wl_r<450> a_wl_r<449> a_wl_r<448>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<59> a_wi<447> a_wi<446> a_wi<445> a_wi<444> a_wi<443> a_wi<442> a_wi<441> a_wi<440> a_wi<439> a_wi<438> a_wi<437> a_wi<436> a_wi<435> a_wi<434> a_wi<433> a_wi<432> a_wl_r<447> a_wl_r<446> a_wl_r<445> a_wl_r<444> a_wl_r<443> a_wl_r<442> a_wl_r<441> a_wl_r<440> a_wl_r<439> a_wl_r<438> a_wl_r<437> a_wl_r<436> a_wl_r<435> a_wl_r<434> a_wl_r<433> a_wl_r<432>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<58> a_wi<431> a_wi<430> a_wi<429> a_wi<428> a_wi<427> a_wi<426> a_wi<425> a_wi<424> a_wi<423> a_wi<422> a_wi<421> a_wi<420> a_wi<419> a_wi<418> a_wi<417> a_wi<416> a_wl_r<431> a_wl_r<430> a_wl_r<429> a_wl_r<428> a_wl_r<427> a_wl_r<426> a_wl_r<425> a_wl_r<424> a_wl_r<423> a_wl_r<422> a_wl_r<421> a_wl_r<420> a_wl_r<419> a_wl_r<418> a_wl_r<417> a_wl_r<416>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<57> a_wi<415> a_wi<414> a_wi<413> a_wi<412> a_wi<411> a_wi<410> a_wi<409> a_wi<408> a_wi<407> a_wi<406> a_wi<405> a_wi<404> a_wi<403> a_wi<402> a_wi<401> a_wi<400> a_wl_r<415> a_wl_r<414> a_wl_r<413> a_wl_r<412> a_wl_r<411> a_wl_r<410> a_wl_r<409> a_wl_r<408> a_wl_r<407> a_wl_r<406> a_wl_r<405> a_wl_r<404> a_wl_r<403> a_wl_r<402> a_wl_r<401> a_wl_r<400>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<56> a_wi<399> a_wi<398> a_wi<397> a_wi<396> a_wi<395> a_wi<394> a_wi<393> a_wi<392> a_wi<391> a_wi<390> a_wi<389> a_wi<388> a_wi<387> a_wi<386> a_wi<385> a_wi<384> a_wl_r<399> a_wl_r<398> a_wl_r<397> a_wl_r<396> a_wl_r<395> a_wl_r<394> a_wl_r<393> a_wl_r<392> a_wl_r<391> a_wl_r<390> a_wl_r<389> a_wl_r<388> a_wl_r<387> a_wl_r<386> a_wl_r<385> a_wl_r<384>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<55> a_wi<383> a_wi<382> a_wi<381> a_wi<380> a_wi<379> a_wi<378> a_wi<377> a_wi<376> a_wi<375> a_wi<374> a_wi<373> a_wi<372> a_wi<371> a_wi<370> a_wi<369> a_wi<368> a_wl_r<383> a_wl_r<382> a_wl_r<381> a_wl_r<380> a_wl_r<379> a_wl_r<378> a_wl_r<377> a_wl_r<376> a_wl_r<375> a_wl_r<374> a_wl_r<373> a_wl_r<372> a_wl_r<371> a_wl_r<370> a_wl_r<369> a_wl_r<368>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<54> a_wi<367> a_wi<366> a_wi<365> a_wi<364> a_wi<363> a_wi<362> a_wi<361> a_wi<360> a_wi<359> a_wi<358> a_wi<357> a_wi<356> a_wi<355> a_wi<354> a_wi<353> a_wi<352> a_wl_r<367> a_wl_r<366> a_wl_r<365> a_wl_r<364> a_wl_r<363> a_wl_r<362> a_wl_r<361> a_wl_r<360> a_wl_r<359> a_wl_r<358> a_wl_r<357> a_wl_r<356> a_wl_r<355> a_wl_r<354> a_wl_r<353> a_wl_r<352>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<53> a_wi<351> a_wi<350> a_wi<349> a_wi<348> a_wi<347> a_wi<346> a_wi<345> a_wi<344> a_wi<343> a_wi<342> a_wi<341> a_wi<340> a_wi<339> a_wi<338> a_wi<337> a_wi<336> a_wl_r<351> a_wl_r<350> a_wl_r<349> a_wl_r<348> a_wl_r<347> a_wl_r<346> a_wl_r<345> a_wl_r<344> a_wl_r<343> a_wl_r<342> a_wl_r<341> a_wl_r<340> a_wl_r<339> a_wl_r<338> a_wl_r<337> a_wl_r<336>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<52> a_wi<335> a_wi<334> a_wi<333> a_wi<332> a_wi<331> a_wi<330> a_wi<329> a_wi<328> a_wi<327> a_wi<326> a_wi<325> a_wi<324> a_wi<323> a_wi<322> a_wi<321> a_wi<320> a_wl_r<335> a_wl_r<334> a_wl_r<333> a_wl_r<332> a_wl_r<331> a_wl_r<330> a_wl_r<329> a_wl_r<328> a_wl_r<327> a_wl_r<326> a_wl_r<325> a_wl_r<324> a_wl_r<323> a_wl_r<322> a_wl_r<321> a_wl_r<320>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<51> a_wi<319> a_wi<318> a_wi<317> a_wi<316> a_wi<315> a_wi<314> a_wi<313> a_wi<312> a_wi<311> a_wi<310> a_wi<309> a_wi<308> a_wi<307> a_wi<306> a_wi<305> a_wi<304> a_wl_r<319> a_wl_r<318> a_wl_r<317> a_wl_r<316> a_wl_r<315> a_wl_r<314> a_wl_r<313> a_wl_r<312> a_wl_r<311> a_wl_r<310> a_wl_r<309> a_wl_r<308> a_wl_r<307> a_wl_r<306> a_wl_r<305> a_wl_r<304>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<50> a_wi<303> a_wi<302> a_wi<301> a_wi<300> a_wi<299> a_wi<298> a_wi<297> a_wi<296> a_wi<295> a_wi<294> a_wi<293> a_wi<292> a_wi<291> a_wi<290> a_wi<289> a_wi<288> a_wl_r<303> a_wl_r<302> a_wl_r<301> a_wl_r<300> a_wl_r<299> a_wl_r<298> a_wl_r<297> a_wl_r<296> a_wl_r<295> a_wl_r<294> a_wl_r<293> a_wl_r<292> a_wl_r<291> a_wl_r<290> a_wl_r<289> a_wl_r<288>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<49> a_wi<287> a_wi<286> a_wi<285> a_wi<284> a_wi<283> a_wi<282> a_wi<281> a_wi<280> a_wi<279> a_wi<278> a_wi<277> a_wi<276> a_wi<275> a_wi<274> a_wi<273> a_wi<272> a_wl_r<287> a_wl_r<286> a_wl_r<285> a_wl_r<284> a_wl_r<283> a_wl_r<282> a_wl_r<281> a_wl_r<280> a_wl_r<279> a_wl_r<278> a_wl_r<277> a_wl_r<276> a_wl_r<275> a_wl_r<274> a_wl_r<273> a_wl_r<272>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<48> a_wi<271> a_wi<270> a_wi<269> a_wi<268> a_wi<267> a_wi<266> a_wi<265> a_wi<264> a_wi<263> a_wi<262> a_wi<261> a_wi<260> a_wi<259> a_wi<258> a_wi<257> a_wi<256> a_wl_r<271> a_wl_r<270> a_wl_r<269> a_wl_r<268> a_wl_r<267> a_wl_r<266> a_wl_r<265> a_wl_r<264> a_wl_r<263> a_wl_r<262> a_wl_r<261> a_wl_r<260> a_wl_r<259> a_wl_r<258> a_wl_r<257> a_wl_r<256>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<47> a_wi<255> a_wi<254> a_wi<253> a_wi<252> a_wi<251> a_wi<250> a_wi<249> a_wi<248> a_wi<247> a_wi<246> a_wi<245> a_wi<244> a_wi<243> a_wi<242> a_wi<241> a_wi<240> a_wl_r<255> a_wl_r<254> a_wl_r<253> a_wl_r<252> a_wl_r<251> a_wl_r<250> a_wl_r<249> a_wl_r<248> a_wl_r<247> a_wl_r<246> a_wl_r<245> a_wl_r<244> a_wl_r<243> a_wl_r<242> a_wl_r<241> a_wl_r<240>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<46> a_wi<239> a_wi<238> a_wi<237> a_wi<236> a_wi<235> a_wi<234> a_wi<233> a_wi<232> a_wi<231> a_wi<230> a_wi<229> a_wi<228> a_wi<227> a_wi<226> a_wi<225> a_wi<224> a_wl_r<239> a_wl_r<238> a_wl_r<237> a_wl_r<236> a_wl_r<235> a_wl_r<234> a_wl_r<233> a_wl_r<232> a_wl_r<231> a_wl_r<230> a_wl_r<229> a_wl_r<228> a_wl_r<227> a_wl_r<226> a_wl_r<225> a_wl_r<224>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<45> a_wi<223> a_wi<222> a_wi<221> a_wi<220> a_wi<219> a_wi<218> a_wi<217> a_wi<216> a_wi<215> a_wi<214> a_wi<213> a_wi<212> a_wi<211> a_wi<210> a_wi<209> a_wi<208> a_wl_r<223> a_wl_r<222> a_wl_r<221> a_wl_r<220> a_wl_r<219> a_wl_r<218> a_wl_r<217> a_wl_r<216> a_wl_r<215> a_wl_r<214> a_wl_r<213> a_wl_r<212> a_wl_r<211> a_wl_r<210> a_wl_r<209> a_wl_r<208>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<44> a_wi<207> a_wi<206> a_wi<205> a_wi<204> a_wi<203> a_wi<202> a_wi<201> a_wi<200> a_wi<199> a_wi<198> a_wi<197> a_wi<196> a_wi<195> a_wi<194> a_wi<193> a_wi<192> a_wl_r<207> a_wl_r<206> a_wl_r<205> a_wl_r<204> a_wl_r<203> a_wl_r<202> a_wl_r<201> a_wl_r<200> a_wl_r<199> a_wl_r<198> a_wl_r<197> a_wl_r<196> a_wl_r<195> a_wl_r<194> a_wl_r<193> a_wl_r<192>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<43> a_wi<191> a_wi<190> a_wi<189> a_wi<188> a_wi<187> a_wi<186> a_wi<185> a_wi<184> a_wi<183> a_wi<182> a_wi<181> a_wi<180> a_wi<179> a_wi<178> a_wi<177> a_wi<176> a_wl_r<191> a_wl_r<190> a_wl_r<189> a_wl_r<188> a_wl_r<187> a_wl_r<186> a_wl_r<185> a_wl_r<184> a_wl_r<183> a_wl_r<182> a_wl_r<181> a_wl_r<180> a_wl_r<179> a_wl_r<178> a_wl_r<177> a_wl_r<176>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<42> a_wi<175> a_wi<174> a_wi<173> a_wi<172> a_wi<171> a_wi<170> a_wi<169> a_wi<168> a_wi<167> a_wi<166> a_wi<165> a_wi<164> a_wi<163> a_wi<162> a_wi<161> a_wi<160> a_wl_r<175> a_wl_r<174> a_wl_r<173> a_wl_r<172> a_wl_r<171> a_wl_r<170> a_wl_r<169> a_wl_r<168> a_wl_r<167> a_wl_r<166> a_wl_r<165> a_wl_r<164> a_wl_r<163> a_wl_r<162> a_wl_r<161> a_wl_r<160>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<41> a_wi<159> a_wi<158> a_wi<157> a_wi<156> a_wi<155> a_wi<154> a_wi<153> a_wi<152> a_wi<151> a_wi<150> a_wi<149> a_wi<148> a_wi<147> a_wi<146> a_wi<145> a_wi<144> a_wl_r<159> a_wl_r<158> a_wl_r<157> a_wl_r<156> a_wl_r<155> a_wl_r<154> a_wl_r<153> a_wl_r<152> a_wl_r<151> a_wl_r<150> a_wl_r<149> a_wl_r<148> a_wl_r<147> a_wl_r<146> a_wl_r<145> a_wl_r<144>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<40> a_wi<143> a_wi<142> a_wi<141> a_wi<140> a_wi<139> a_wi<138> a_wi<137> a_wi<136> a_wi<135> a_wi<134> a_wi<133> a_wi<132> a_wi<131> a_wi<130> a_wi<129> a_wi<128> a_wl_r<143> a_wl_r<142> a_wl_r<141> a_wl_r<140> a_wl_r<139> a_wl_r<138> a_wl_r<137> a_wl_r<136> a_wl_r<135> a_wl_r<134> a_wl_r<133> a_wl_r<132> a_wl_r<131> a_wl_r<130> a_wl_r<129> a_wl_r<128>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<39> a_wi<127> a_wi<126> a_wi<125> a_wi<124> a_wi<123> a_wi<122> a_wi<121> a_wi<120> a_wi<119> a_wi<118> a_wi<117> a_wi<116> a_wi<115> a_wi<114> a_wi<113> a_wi<112> a_wl_r<127> a_wl_r<126> a_wl_r<125> a_wl_r<124> a_wl_r<123> a_wl_r<122> a_wl_r<121> a_wl_r<120> a_wl_r<119> a_wl_r<118> a_wl_r<117> a_wl_r<116> a_wl_r<115> a_wl_r<114> a_wl_r<113> a_wl_r<112>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<38> a_wi<111> a_wi<110> a_wi<109> a_wi<108> a_wi<107> a_wi<106> a_wi<105> a_wi<104> a_wi<103> a_wi<102> a_wi<101> a_wi<100> a_wi<99> a_wi<98> a_wi<97> a_wi<96> a_wl_r<111> a_wl_r<110> a_wl_r<109> a_wl_r<108> a_wl_r<107> a_wl_r<106> a_wl_r<105> a_wl_r<104> a_wl_r<103> a_wl_r<102> a_wl_r<101> a_wl_r<100> a_wl_r<99> a_wl_r<98> a_wl_r<97> a_wl_r<96>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<37> a_wi<95> a_wi<94> a_wi<93> a_wi<92> a_wi<91> a_wi<90> a_wi<89> a_wi<88> a_wi<87> a_wi<86> a_wi<85> a_wi<84> a_wi<83> a_wi<82> a_wi<81> a_wi<80> a_wl_r<95> a_wl_r<94> a_wl_r<93> a_wl_r<92> a_wl_r<91> a_wl_r<90> a_wl_r<89> a_wl_r<88> a_wl_r<87> a_wl_r<86> a_wl_r<85> a_wl_r<84> a_wl_r<83> a_wl_r<82> a_wl_r<81> a_wl_r<80>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<36> a_wi<79> a_wi<78> a_wi<77> a_wi<76> a_wi<75> a_wi<74> a_wi<73> a_wi<72> a_wi<71> a_wi<70> a_wi<69> a_wi<68> a_wi<67> a_wi<66> a_wi<65> a_wi<64> a_wl_r<79> a_wl_r<78> a_wl_r<77> a_wl_r<76> a_wl_r<75> a_wl_r<74> a_wl_r<73> a_wl_r<72> a_wl_r<71> a_wl_r<70> a_wl_r<69> a_wl_r<68> a_wl_r<67> a_wl_r<66> a_wl_r<65> a_wl_r<64>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<35> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wl_r<63> a_wl_r<62> a_wl_r<61> a_wl_r<60> a_wl_r<59> a_wl_r<58> a_wl_r<57> a_wl_r<56> a_wl_r<55> a_wl_r<54> a_wl_r<53> a_wl_r<52> a_wl_r<51> a_wl_r<50> a_wl_r<49> a_wl_r<48>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<34> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wl_r<47> a_wl_r<46> a_wl_r<45> a_wl_r<44> a_wl_r<43> a_wl_r<42> a_wl_r<41> a_wl_r<40> a_wl_r<39> a_wl_r<38> a_wl_r<37> a_wl_r<36> a_wl_r<35> a_wl_r<34> a_wl_r<33> a_wl_r<32>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<33> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wl_r<31> a_wl_r<30> a_wl_r<29> a_wl_r<28> a_wl_r<27> a_wl_r<26> a_wl_r<25> a_wl_r<24> a_wl_r<23> a_wl_r<22> a_wl_r<21> a_wl_r<20> a_wl_r<19> a_wl_r<18> a_wl_r<17> a_wl_r<16>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<32> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> a_wl_r<15> a_wl_r<14> a_wl_r<13> a_wl_r<12> a_wl_r<11> a_wl_r<10> a_wl_r<9> a_wl_r<8> a_wl_r<7> a_wl_r<6> a_wl_r<5> a_wl_r<4> a_wl_r<3> a_wl_r<2> a_wl_r<1> a_wl_r<0>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<31> a_wi<511> a_wi<510> a_wi<509> a_wi<508> a_wi<507> a_wi<506> a_wi<505> a_wi<504> a_wi<503> a_wi<502> a_wi<501> a_wi<500> a_wi<499> a_wi<498> a_wi<497> a_wi<496> a_wl_l<511> a_wl_l<510> a_wl_l<509> a_wl_l<508> a_wl_l<507> a_wl_l<506> a_wl_l<505> a_wl_l<504> a_wl_l<503> a_wl_l<502> a_wl_l<501> a_wl_l<500> a_wl_l<499> a_wl_l<498> a_wl_l<497> a_wl_l<496>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<30> a_wi<495> a_wi<494> a_wi<493> a_wi<492> a_wi<491> a_wi<490> a_wi<489> a_wi<488> a_wi<487> a_wi<486> a_wi<485> a_wi<484> a_wi<483> a_wi<482> a_wi<481> a_wi<480> a_wl_l<495> a_wl_l<494> a_wl_l<493> a_wl_l<492> a_wl_l<491> a_wl_l<490> a_wl_l<489> a_wl_l<488> a_wl_l<487> a_wl_l<486> a_wl_l<485> a_wl_l<484> a_wl_l<483> a_wl_l<482> a_wl_l<481> a_wl_l<480>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<29> a_wi<479> a_wi<478> a_wi<477> a_wi<476> a_wi<475> a_wi<474> a_wi<473> a_wi<472> a_wi<471> a_wi<470> a_wi<469> a_wi<468> a_wi<467> a_wi<466> a_wi<465> a_wi<464> a_wl_l<479> a_wl_l<478> a_wl_l<477> a_wl_l<476> a_wl_l<475> a_wl_l<474> a_wl_l<473> a_wl_l<472> a_wl_l<471> a_wl_l<470> a_wl_l<469> a_wl_l<468> a_wl_l<467> a_wl_l<466> a_wl_l<465> a_wl_l<464>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<28> a_wi<463> a_wi<462> a_wi<461> a_wi<460> a_wi<459> a_wi<458> a_wi<457> a_wi<456> a_wi<455> a_wi<454> a_wi<453> a_wi<452> a_wi<451> a_wi<450> a_wi<449> a_wi<448> a_wl_l<463> a_wl_l<462> a_wl_l<461> a_wl_l<460> a_wl_l<459> a_wl_l<458> a_wl_l<457> a_wl_l<456> a_wl_l<455> a_wl_l<454> a_wl_l<453> a_wl_l<452> a_wl_l<451> a_wl_l<450> a_wl_l<449> a_wl_l<448>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<27> a_wi<447> a_wi<446> a_wi<445> a_wi<444> a_wi<443> a_wi<442> a_wi<441> a_wi<440> a_wi<439> a_wi<438> a_wi<437> a_wi<436> a_wi<435> a_wi<434> a_wi<433> a_wi<432> a_wl_l<447> a_wl_l<446> a_wl_l<445> a_wl_l<444> a_wl_l<443> a_wl_l<442> a_wl_l<441> a_wl_l<440> a_wl_l<439> a_wl_l<438> a_wl_l<437> a_wl_l<436> a_wl_l<435> a_wl_l<434> a_wl_l<433> a_wl_l<432>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<26> a_wi<431> a_wi<430> a_wi<429> a_wi<428> a_wi<427> a_wi<426> a_wi<425> a_wi<424> a_wi<423> a_wi<422> a_wi<421> a_wi<420> a_wi<419> a_wi<418> a_wi<417> a_wi<416> a_wl_l<431> a_wl_l<430> a_wl_l<429> a_wl_l<428> a_wl_l<427> a_wl_l<426> a_wl_l<425> a_wl_l<424> a_wl_l<423> a_wl_l<422> a_wl_l<421> a_wl_l<420> a_wl_l<419> a_wl_l<418> a_wl_l<417> a_wl_l<416>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<25> a_wi<415> a_wi<414> a_wi<413> a_wi<412> a_wi<411> a_wi<410> a_wi<409> a_wi<408> a_wi<407> a_wi<406> a_wi<405> a_wi<404> a_wi<403> a_wi<402> a_wi<401> a_wi<400> a_wl_l<415> a_wl_l<414> a_wl_l<413> a_wl_l<412> a_wl_l<411> a_wl_l<410> a_wl_l<409> a_wl_l<408> a_wl_l<407> a_wl_l<406> a_wl_l<405> a_wl_l<404> a_wl_l<403> a_wl_l<402> a_wl_l<401> a_wl_l<400>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<24> a_wi<399> a_wi<398> a_wi<397> a_wi<396> a_wi<395> a_wi<394> a_wi<393> a_wi<392> a_wi<391> a_wi<390> a_wi<389> a_wi<388> a_wi<387> a_wi<386> a_wi<385> a_wi<384> a_wl_l<399> a_wl_l<398> a_wl_l<397> a_wl_l<396> a_wl_l<395> a_wl_l<394> a_wl_l<393> a_wl_l<392> a_wl_l<391> a_wl_l<390> a_wl_l<389> a_wl_l<388> a_wl_l<387> a_wl_l<386> a_wl_l<385> a_wl_l<384>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<23> a_wi<383> a_wi<382> a_wi<381> a_wi<380> a_wi<379> a_wi<378> a_wi<377> a_wi<376> a_wi<375> a_wi<374> a_wi<373> a_wi<372> a_wi<371> a_wi<370> a_wi<369> a_wi<368> a_wl_l<383> a_wl_l<382> a_wl_l<381> a_wl_l<380> a_wl_l<379> a_wl_l<378> a_wl_l<377> a_wl_l<376> a_wl_l<375> a_wl_l<374> a_wl_l<373> a_wl_l<372> a_wl_l<371> a_wl_l<370> a_wl_l<369> a_wl_l<368>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<22> a_wi<367> a_wi<366> a_wi<365> a_wi<364> a_wi<363> a_wi<362> a_wi<361> a_wi<360> a_wi<359> a_wi<358> a_wi<357> a_wi<356> a_wi<355> a_wi<354> a_wi<353> a_wi<352> a_wl_l<367> a_wl_l<366> a_wl_l<365> a_wl_l<364> a_wl_l<363> a_wl_l<362> a_wl_l<361> a_wl_l<360> a_wl_l<359> a_wl_l<358> a_wl_l<357> a_wl_l<356> a_wl_l<355> a_wl_l<354> a_wl_l<353> a_wl_l<352>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<21> a_wi<351> a_wi<350> a_wi<349> a_wi<348> a_wi<347> a_wi<346> a_wi<345> a_wi<344> a_wi<343> a_wi<342> a_wi<341> a_wi<340> a_wi<339> a_wi<338> a_wi<337> a_wi<336> a_wl_l<351> a_wl_l<350> a_wl_l<349> a_wl_l<348> a_wl_l<347> a_wl_l<346> a_wl_l<345> a_wl_l<344> a_wl_l<343> a_wl_l<342> a_wl_l<341> a_wl_l<340> a_wl_l<339> a_wl_l<338> a_wl_l<337> a_wl_l<336>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<20> a_wi<335> a_wi<334> a_wi<333> a_wi<332> a_wi<331> a_wi<330> a_wi<329> a_wi<328> a_wi<327> a_wi<326> a_wi<325> a_wi<324> a_wi<323> a_wi<322> a_wi<321> a_wi<320> a_wl_l<335> a_wl_l<334> a_wl_l<333> a_wl_l<332> a_wl_l<331> a_wl_l<330> a_wl_l<329> a_wl_l<328> a_wl_l<327> a_wl_l<326> a_wl_l<325> a_wl_l<324> a_wl_l<323> a_wl_l<322> a_wl_l<321> a_wl_l<320>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<19> a_wi<319> a_wi<318> a_wi<317> a_wi<316> a_wi<315> a_wi<314> a_wi<313> a_wi<312> a_wi<311> a_wi<310> a_wi<309> a_wi<308> a_wi<307> a_wi<306> a_wi<305> a_wi<304> a_wl_l<319> a_wl_l<318> a_wl_l<317> a_wl_l<316> a_wl_l<315> a_wl_l<314> a_wl_l<313> a_wl_l<312> a_wl_l<311> a_wl_l<310> a_wl_l<309> a_wl_l<308> a_wl_l<307> a_wl_l<306> a_wl_l<305> a_wl_l<304>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<18> a_wi<303> a_wi<302> a_wi<301> a_wi<300> a_wi<299> a_wi<298> a_wi<297> a_wi<296> a_wi<295> a_wi<294> a_wi<293> a_wi<292> a_wi<291> a_wi<290> a_wi<289> a_wi<288> a_wl_l<303> a_wl_l<302> a_wl_l<301> a_wl_l<300> a_wl_l<299> a_wl_l<298> a_wl_l<297> a_wl_l<296> a_wl_l<295> a_wl_l<294> a_wl_l<293> a_wl_l<292> a_wl_l<291> a_wl_l<290> a_wl_l<289> a_wl_l<288>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<17> a_wi<287> a_wi<286> a_wi<285> a_wi<284> a_wi<283> a_wi<282> a_wi<281> a_wi<280> a_wi<279> a_wi<278> a_wi<277> a_wi<276> a_wi<275> a_wi<274> a_wi<273> a_wi<272> a_wl_l<287> a_wl_l<286> a_wl_l<285> a_wl_l<284> a_wl_l<283> a_wl_l<282> a_wl_l<281> a_wl_l<280> a_wl_l<279> a_wl_l<278> a_wl_l<277> a_wl_l<276> a_wl_l<275> a_wl_l<274> a_wl_l<273> a_wl_l<272>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<16> a_wi<271> a_wi<270> a_wi<269> a_wi<268> a_wi<267> a_wi<266> a_wi<265> a_wi<264> a_wi<263> a_wi<262> a_wi<261> a_wi<260> a_wi<259> a_wi<258> a_wi<257> a_wi<256> a_wl_l<271> a_wl_l<270> a_wl_l<269> a_wl_l<268> a_wl_l<267> a_wl_l<266> a_wl_l<265> a_wl_l<264> a_wl_l<263> a_wl_l<262> a_wl_l<261> a_wl_l<260> a_wl_l<259> a_wl_l<258> a_wl_l<257> a_wl_l<256>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<15> a_wi<255> a_wi<254> a_wi<253> a_wi<252> a_wi<251> a_wi<250> a_wi<249> a_wi<248> a_wi<247> a_wi<246> a_wi<245> a_wi<244> a_wi<243> a_wi<242> a_wi<241> a_wi<240> a_wl_l<255> a_wl_l<254> a_wl_l<253> a_wl_l<252> a_wl_l<251> a_wl_l<250> a_wl_l<249> a_wl_l<248> a_wl_l<247> a_wl_l<246> a_wl_l<245> a_wl_l<244> a_wl_l<243> a_wl_l<242> a_wl_l<241> a_wl_l<240>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<14> a_wi<239> a_wi<238> a_wi<237> a_wi<236> a_wi<235> a_wi<234> a_wi<233> a_wi<232> a_wi<231> a_wi<230> a_wi<229> a_wi<228> a_wi<227> a_wi<226> a_wi<225> a_wi<224> a_wl_l<239> a_wl_l<238> a_wl_l<237> a_wl_l<236> a_wl_l<235> a_wl_l<234> a_wl_l<233> a_wl_l<232> a_wl_l<231> a_wl_l<230> a_wl_l<229> a_wl_l<228> a_wl_l<227> a_wl_l<226> a_wl_l<225> a_wl_l<224>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<13> a_wi<223> a_wi<222> a_wi<221> a_wi<220> a_wi<219> a_wi<218> a_wi<217> a_wi<216> a_wi<215> a_wi<214> a_wi<213> a_wi<212> a_wi<211> a_wi<210> a_wi<209> a_wi<208> a_wl_l<223> a_wl_l<222> a_wl_l<221> a_wl_l<220> a_wl_l<219> a_wl_l<218> a_wl_l<217> a_wl_l<216> a_wl_l<215> a_wl_l<214> a_wl_l<213> a_wl_l<212> a_wl_l<211> a_wl_l<210> a_wl_l<209> a_wl_l<208>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<12> a_wi<207> a_wi<206> a_wi<205> a_wi<204> a_wi<203> a_wi<202> a_wi<201> a_wi<200> a_wi<199> a_wi<198> a_wi<197> a_wi<196> a_wi<195> a_wi<194> a_wi<193> a_wi<192> a_wl_l<207> a_wl_l<206> a_wl_l<205> a_wl_l<204> a_wl_l<203> a_wl_l<202> a_wl_l<201> a_wl_l<200> a_wl_l<199> a_wl_l<198> a_wl_l<197> a_wl_l<196> a_wl_l<195> a_wl_l<194> a_wl_l<193> a_wl_l<192>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<11> a_wi<191> a_wi<190> a_wi<189> a_wi<188> a_wi<187> a_wi<186> a_wi<185> a_wi<184> a_wi<183> a_wi<182> a_wi<181> a_wi<180> a_wi<179> a_wi<178> a_wi<177> a_wi<176> a_wl_l<191> a_wl_l<190> a_wl_l<189> a_wl_l<188> a_wl_l<187> a_wl_l<186> a_wl_l<185> a_wl_l<184> a_wl_l<183> a_wl_l<182> a_wl_l<181> a_wl_l<180> a_wl_l<179> a_wl_l<178> a_wl_l<177> a_wl_l<176>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<10> a_wi<175> a_wi<174> a_wi<173> a_wi<172> a_wi<171> a_wi<170> a_wi<169> a_wi<168> a_wi<167> a_wi<166> a_wi<165> a_wi<164> a_wi<163> a_wi<162> a_wi<161> a_wi<160> a_wl_l<175> a_wl_l<174> a_wl_l<173> a_wl_l<172> a_wl_l<171> a_wl_l<170> a_wl_l<169> a_wl_l<168> a_wl_l<167> a_wl_l<166> a_wl_l<165> a_wl_l<164> a_wl_l<163> a_wl_l<162> a_wl_l<161> a_wl_l<160>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<9> a_wi<159> a_wi<158> a_wi<157> a_wi<156> a_wi<155> a_wi<154> a_wi<153> a_wi<152> a_wi<151> a_wi<150> a_wi<149> a_wi<148> a_wi<147> a_wi<146> a_wi<145> a_wi<144> a_wl_l<159> a_wl_l<158> a_wl_l<157> a_wl_l<156> a_wl_l<155> a_wl_l<154> a_wl_l<153> a_wl_l<152> a_wl_l<151> a_wl_l<150> a_wl_l<149> a_wl_l<148> a_wl_l<147> a_wl_l<146> a_wl_l<145> a_wl_l<144>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<8> a_wi<143> a_wi<142> a_wi<141> a_wi<140> a_wi<139> a_wi<138> a_wi<137> a_wi<136> a_wi<135> a_wi<134> a_wi<133> a_wi<132> a_wi<131> a_wi<130> a_wi<129> a_wi<128> a_wl_l<143> a_wl_l<142> a_wl_l<141> a_wl_l<140> a_wl_l<139> a_wl_l<138> a_wl_l<137> a_wl_l<136> a_wl_l<135> a_wl_l<134> a_wl_l<133> a_wl_l<132> a_wl_l<131> a_wl_l<130> a_wl_l<129> a_wl_l<128>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<7> a_wi<127> a_wi<126> a_wi<125> a_wi<124> a_wi<123> a_wi<122> a_wi<121> a_wi<120> a_wi<119> a_wi<118> a_wi<117> a_wi<116> a_wi<115> a_wi<114> a_wi<113> a_wi<112> a_wl_l<127> a_wl_l<126> a_wl_l<125> a_wl_l<124> a_wl_l<123> a_wl_l<122> a_wl_l<121> a_wl_l<120> a_wl_l<119> a_wl_l<118> a_wl_l<117> a_wl_l<116> a_wl_l<115> a_wl_l<114> a_wl_l<113> a_wl_l<112>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<6> a_wi<111> a_wi<110> a_wi<109> a_wi<108> a_wi<107> a_wi<106> a_wi<105> a_wi<104> a_wi<103> a_wi<102> a_wi<101> a_wi<100> a_wi<99> a_wi<98> a_wi<97> a_wi<96> a_wl_l<111> a_wl_l<110> a_wl_l<109> a_wl_l<108> a_wl_l<107> a_wl_l<106> a_wl_l<105> a_wl_l<104> a_wl_l<103> a_wl_l<102> a_wl_l<101> a_wl_l<100> a_wl_l<99> a_wl_l<98> a_wl_l<97> a_wl_l<96>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<5> a_wi<95> a_wi<94> a_wi<93> a_wi<92> a_wi<91> a_wi<90> a_wi<89> a_wi<88> a_wi<87> a_wi<86> a_wi<85> a_wi<84> a_wi<83> a_wi<82> a_wi<81> a_wi<80> a_wl_l<95> a_wl_l<94> a_wl_l<93> a_wl_l<92> a_wl_l<91> a_wl_l<90> a_wl_l<89> a_wl_l<88> a_wl_l<87> a_wl_l<86> a_wl_l<85> a_wl_l<84> a_wl_l<83> a_wl_l<82> a_wl_l<81> a_wl_l<80>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<4> a_wi<79> a_wi<78> a_wi<77> a_wi<76> a_wi<75> a_wi<74> a_wi<73> a_wi<72> a_wi<71> a_wi<70> a_wi<69> a_wi<68> a_wi<67> a_wi<66> a_wi<65> a_wi<64> a_wl_l<79> a_wl_l<78> a_wl_l<77> a_wl_l<76> a_wl_l<75> a_wl_l<74> a_wl_l<73> a_wl_l<72> a_wl_l<71> a_wl_l<70> a_wl_l<69> a_wl_l<68> a_wl_l<67> a_wl_l<66> a_wl_l<65> a_wl_l<64>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<3> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wl_l<63> a_wl_l<62> a_wl_l<61> a_wl_l<60> a_wl_l<59> a_wl_l<58> a_wl_l<57> a_wl_l<56> a_wl_l<55> a_wl_l<54> a_wl_l<53> a_wl_l<52> a_wl_l<51> a_wl_l<50> a_wl_l<49> a_wl_l<48>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<2> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wl_l<47> a_wl_l<46> a_wl_l<45> a_wl_l<44> a_wl_l<43> a_wl_l<42> a_wl_l<41> a_wl_l<40> a_wl_l<39> a_wl_l<38> a_wl_l<37> a_wl_l<36> a_wl_l<35> a_wl_l<34> a_wl_l<33> a_wl_l<32>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<1> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wl_l<31> a_wl_l<30> a_wl_l<29> a_wl_l<28> a_wl_l<27> a_wl_l<26> a_wl_l<25> a_wl_l<24> a_wl_l<23> a_wl_l<22> a_wl_l<21> a_wl_l<20> a_wl_l<19> a_wl_l<18> a_wl_l<17> a_wl_l<16>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8
XA_WLDRV<0> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> a_wl_l<15> a_wl_l<14> a_wl_l<13> a_wl_l<12> a_wl_l<11> a_wl_l<10> a_wl_l<9> a_wl_l<8> a_wl_l<7> a_wl_l<6> a_wl_l<5> a_wl_l<4> a_wl_l<3> a_wl_l<2> a_wl_l<1> a_wl_l<0>  VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_WLDRV16X8


XA_CTRL a_aclk_n A_BIST_CLK A_BIST_MEN A_BIST_EN A_BIST_REN A_BIST_WEN a_tiel A_CLK A_MEN a_dclk a_eclk a_pulse_h a_pulse_l a_pulse a_rclk A_REN a_cs a_wclk A_WEN VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_CTRL


XA_ROWDEC a_addr_row<8> a_addr_row<7> a_addr_row<6> a_addr_row<5> a_addr_row<4> a_addr_row<3> a_addr_row<2> a_addr_row<1> a_addr_row<0> a_cs a_eclk a_wi<511> a_wi<510> a_wi<509> a_wi<508> a_wi<507> a_wi<506> a_wi<505> a_wi<504> a_wi<503> a_wi<502> a_wi<501> a_wi<500> a_wi<499> a_wi<498> a_wi<497> a_wi<496> a_wi<495> a_wi<494> a_wi<493> a_wi<492> a_wi<491> a_wi<490> a_wi<489> a_wi<488> a_wi<487> a_wi<486> a_wi<485> a_wi<484> a_wi<483> a_wi<482> a_wi<481> a_wi<480> a_wi<479> a_wi<478> a_wi<477> a_wi<476> a_wi<475> a_wi<474> a_wi<473> a_wi<472> a_wi<471> a_wi<470> a_wi<469> a_wi<468> a_wi<467> a_wi<466> a_wi<465> a_wi<464> a_wi<463> a_wi<462> a_wi<461> a_wi<460> a_wi<459> a_wi<458> a_wi<457> a_wi<456> a_wi<455> a_wi<454> a_wi<453> a_wi<452> a_wi<451> a_wi<450> a_wi<449> a_wi<448> a_wi<447> a_wi<446> a_wi<445> a_wi<444> a_wi<443> a_wi<442> a_wi<441> a_wi<440> a_wi<439> a_wi<438> a_wi<437> a_wi<436> a_wi<435> a_wi<434> a_wi<433> a_wi<432> a_wi<431> a_wi<430> a_wi<429> a_wi<428> a_wi<427> a_wi<426> a_wi<425> a_wi<424> a_wi<423> a_wi<422> a_wi<421> a_wi<420> a_wi<419> a_wi<418> a_wi<417> a_wi<416> a_wi<415> a_wi<414> a_wi<413> a_wi<412> a_wi<411> a_wi<410> a_wi<409> a_wi<408> a_wi<407> a_wi<406> a_wi<405> a_wi<404> a_wi<403> a_wi<402> a_wi<401> a_wi<400> a_wi<399> a_wi<398> a_wi<397> a_wi<396> a_wi<395> a_wi<394> a_wi<393> a_wi<392> a_wi<391> a_wi<390> a_wi<389> a_wi<388> a_wi<387> a_wi<386> a_wi<385> a_wi<384> a_wi<383> a_wi<382> a_wi<381> a_wi<380> a_wi<379> a_wi<378> a_wi<377> a_wi<376> a_wi<375> a_wi<374> a_wi<373> a_wi<372> a_wi<371> a_wi<370> a_wi<369> a_wi<368> a_wi<367> a_wi<366> a_wi<365> a_wi<364> a_wi<363> a_wi<362> a_wi<361> a_wi<360> a_wi<359> a_wi<358> a_wi<357> a_wi<356> a_wi<355> a_wi<354> a_wi<353> a_wi<352> a_wi<351> a_wi<350> a_wi<349> a_wi<348> a_wi<347> a_wi<346> a_wi<345> a_wi<344> a_wi<343> a_wi<342> a_wi<341> a_wi<340> a_wi<339> a_wi<338> a_wi<337> a_wi<336> a_wi<335> a_wi<334> a_wi<333> a_wi<332> a_wi<331> a_wi<330> a_wi<329> a_wi<328> a_wi<327> a_wi<326> a_wi<325> a_wi<324> a_wi<323> a_wi<322> a_wi<321> a_wi<320> a_wi<319> a_wi<318> a_wi<317> a_wi<316> a_wi<315> a_wi<314> a_wi<313> a_wi<312> a_wi<311> a_wi<310> a_wi<309> a_wi<308> a_wi<307> a_wi<306> a_wi<305> a_wi<304> a_wi<303> a_wi<302> a_wi<301> a_wi<300> a_wi<299> a_wi<298> a_wi<297> a_wi<296> a_wi<295> a_wi<294> a_wi<293> a_wi<292> a_wi<291> a_wi<290> a_wi<289> a_wi<288> a_wi<287> a_wi<286> a_wi<285> a_wi<284> a_wi<283> a_wi<282> a_wi<281> a_wi<280> a_wi<279> a_wi<278> a_wi<277> a_wi<276> a_wi<275> a_wi<274> a_wi<273> a_wi<272> a_wi<271> a_wi<270> a_wi<269> a_wi<268> a_wi<267> a_wi<266> a_wi<265> a_wi<264> a_wi<263> a_wi<262> a_wi<261> a_wi<260> a_wi<259> a_wi<258> a_wi<257> a_wi<256> a_wi<255> a_wi<254> a_wi<253> a_wi<252> a_wi<251> a_wi<250> a_wi<249> a_wi<248> a_wi<247> a_wi<246> a_wi<245> a_wi<244> a_wi<243> a_wi<242> a_wi<241> a_wi<240> a_wi<239> a_wi<238> a_wi<237> a_wi<236> a_wi<235> a_wi<234> a_wi<233> a_wi<232> a_wi<231> a_wi<230> a_wi<229> a_wi<228> a_wi<227> a_wi<226> a_wi<225> a_wi<224> a_wi<223> a_wi<222> a_wi<221> a_wi<220> a_wi<219> a_wi<218> a_wi<217> a_wi<216> a_wi<215> a_wi<214> a_wi<213> a_wi<212> a_wi<211> a_wi<210> a_wi<209> a_wi<208> a_wi<207> a_wi<206> a_wi<205> a_wi<204> a_wi<203> a_wi<202> a_wi<201> a_wi<200> a_wi<199> a_wi<198> a_wi<197> a_wi<196> a_wi<195> a_wi<194> a_wi<193> a_wi<192> a_wi<191> a_wi<190> a_wi<189> a_wi<188> a_wi<187> a_wi<186> a_wi<185> a_wi<184> a_wi<183> a_wi<182> a_wi<181> a_wi<180> a_wi<179> a_wi<178> a_wi<177> a_wi<176> a_wi<175> a_wi<174> a_wi<173> a_wi<172> a_wi<171> a_wi<170> a_wi<169> a_wi<168> a_wi<167> a_wi<166> a_wi<165> a_wi<164> a_wi<163> a_wi<162> a_wi<161> a_wi<160> a_wi<159> a_wi<158> a_wi<157> a_wi<156> a_wi<155> a_wi<154> a_wi<153> a_wi<152> a_wi<151> a_wi<150> a_wi<149> a_wi<148> a_wi<147> a_wi<146> a_wi<145> a_wi<144> a_wi<143> a_wi<142> a_wi<141> a_wi<140> a_wi<139> a_wi<138> a_wi<137> a_wi<136> a_wi<135> a_wi<134> a_wi<133> a_wi<132> a_wi<131> a_wi<130> a_wi<129> a_wi<128> a_wi<127> a_wi<126> a_wi<125> a_wi<124> a_wi<123> a_wi<122> a_wi<121> a_wi<120> a_wi<119> a_wi<118> a_wi<117> a_wi<116> a_wi<115> a_wi<114> a_wi<113> a_wi<112> a_wi<111> a_wi<110> a_wi<109> a_wi<108> a_wi<107> a_wi<106> a_wi<105> a_wi<104> a_wi<103> a_wi<102> a_wi<101> a_wi<100> a_wi<99> a_wi<98> a_wi<97> a_wi<96> a_wi<95> a_wi<94> a_wi<93> a_wi<92> a_wi<91> a_wi<90> a_wi<89> a_wi<88> a_wi<87> a_wi<86> a_wi<85> a_wi<84> a_wi<83> a_wi<82> a_wi<81> a_wi<80> a_wi<79> a_wi<78> a_wi<77> a_wi<76> a_wi<75> a_wi<74> a_wi<73> a_wi<72> a_wi<71> a_wi<70> a_wi<69> a_wi<68> a_wi<67> a_wi<66> a_wi<65> a_wi<64> a_wi<63> a_wi<62> a_wi<61> a_wi<60> a_wi<59> a_wi<58> a_wi<57> a_wi<56> a_wi<55> a_wi<54> a_wi<53> a_wi<52> a_wi<51> a_wi<50> a_wi<49> a_wi<48> a_wi<47> a_wi<46> a_wi<45> a_wi<44> a_wi<43> a_wi<42> a_wi<41> a_wi<40> a_wi<39> a_wi<38> a_wi<37> a_wi<36> a_wi<35> a_wi<34> a_wi<33> a_wi<32> a_wi<31> a_wi<30> a_wi<29> a_wi<28> a_wi<27> a_wi<26> a_wi<25> a_wi<24> a_wi<23> a_wi<22> a_wi<21> a_wi<20> a_wi<19> a_wi<18> a_wi<17> a_wi<16> a_wi<15> a_wi<14> a_wi<13> a_wi<12> a_wi<11> a_wi<10> a_wi<9> a_wi<8> a_wi<7> a_wi<6> a_wi<5> a_wi<4> a_wi<3> a_wi<2> a_wi<1> a_wi<0> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_ROWDEC9
XA_ROWREG a_aclk_n A_ADDR<10> A_ADDR<9> A_ADDR<8> A_ADDR<7> A_ADDR<6> A_ADDR<5> A_ADDR<4> A_ADDR<3> A_ADDR<2> a_addr_row<8> a_addr_row<7> a_addr_row<6> a_addr_row<5> a_addr_row<4> a_addr_row<3> a_addr_row<2> a_addr_row<1> a_addr_row<0> A_BIST_ADDR<10> A_BIST_ADDR<9> A_BIST_ADDR<8> A_BIST_ADDR<7> A_BIST_ADDR<6> A_BIST_ADDR<5> A_BIST_ADDR<4> A_BIST_ADDR<3> A_BIST_ADDR<2> A_BIST_EN VDD! VSS!  / RM_IHPSG13_2048x64_c2_1P_ROWREG9
XA_COLDEC a_aclk_n A_ADDR<1> A_ADDR<0> a_addr_col<1> a_addr_col<0> a_addr_dec<7> a_addr_dec<6> a_addr_dec<5> a_addr_dec<4> a_addr_dec<3> a_addr_dec<2> a_addr_dec<1> a_addr_dec<0> A_BIST_ADDR<1> A_BIST_ADDR<0> A_BIST_EN VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDEC2


XA_DLYH a_pulse a_pulse_h VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_DLY_pcell_2
XA_DLYL a_pulse_x a_pulse_l VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_DLY_pcell_3
XA_DLYMUX a_pulse_h A_DLY a_pulse_x VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_DLY_MUX

XCOLCTRL<63> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<63> A_BIST_DIN<63> A_BIST_EN a_blc_r<127> a_blc_r<126> a_blc_r<125> a_blc_r<124> a_blt_r<127> a_blt_r<126> a_blt_r<125> a_blt_r<124> A_BM<63> a_dclk_n_r<31> a_dclk_n_r<32> a_dclk_p_r<31> a_dclk_p_r<32> A_DOUT<63> A_DIN<63> a_rclk_n_r<31> a_rclk_n_r<32> a_rclk_p_r<31> a_rclk_p_r<32> a_tieh<63> a_wclk_n_r<31> a_wclk_n_r<32> a_wclk_p_r<31> a_wclk_p_r<32> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<62> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<62> A_BIST_DIN<62> A_BIST_EN a_blc_r<123> a_blc_r<122> a_blc_r<121> a_blc_r<120> a_blt_r<123> a_blt_r<122> a_blt_r<121> a_blt_r<120> A_BM<62> a_dclk_n_r<30> a_dclk_n_r<31> a_dclk_p_r<30> a_dclk_p_r<31> A_DOUT<62> A_DIN<62> a_rclk_n_r<30> a_rclk_n_r<31> a_rclk_p_r<30> a_rclk_p_r<31> a_tieh<62> a_wclk_n_r<30> a_wclk_n_r<31> a_wclk_p_r<30> a_wclk_p_r<31> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<61> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<61> A_BIST_DIN<61> A_BIST_EN a_blc_r<119> a_blc_r<118> a_blc_r<117> a_blc_r<116> a_blt_r<119> a_blt_r<118> a_blt_r<117> a_blt_r<116> A_BM<61> a_dclk_n_r<29> a_dclk_n_r<30> a_dclk_p_r<29> a_dclk_p_r<30> A_DOUT<61> A_DIN<61> a_rclk_n_r<29> a_rclk_n_r<30> a_rclk_p_r<29> a_rclk_p_r<30> a_tieh<61> a_wclk_n_r<29> a_wclk_n_r<30> a_wclk_p_r<29> a_wclk_p_r<30> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<60> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<60> A_BIST_DIN<60> A_BIST_EN a_blc_r<115> a_blc_r<114> a_blc_r<113> a_blc_r<112> a_blt_r<115> a_blt_r<114> a_blt_r<113> a_blt_r<112> A_BM<60> a_dclk_n_r<28> a_dclk_n_r<29> a_dclk_p_r<28> a_dclk_p_r<29> A_DOUT<60> A_DIN<60> a_rclk_n_r<28> a_rclk_n_r<29> a_rclk_p_r<28> a_rclk_p_r<29> a_tieh<60> a_wclk_n_r<28> a_wclk_n_r<29> a_wclk_p_r<28> a_wclk_p_r<29> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<59> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<59> A_BIST_DIN<59> A_BIST_EN a_blc_r<111> a_blc_r<110> a_blc_r<109> a_blc_r<108> a_blt_r<111> a_blt_r<110> a_blt_r<109> a_blt_r<108> A_BM<59> a_dclk_n_r<27> a_dclk_n_r<28> a_dclk_p_r<27> a_dclk_p_r<28> A_DOUT<59> A_DIN<59> a_rclk_n_r<27> a_rclk_n_r<28> a_rclk_p_r<27> a_rclk_p_r<28> a_tieh<59> a_wclk_n_r<27> a_wclk_n_r<28> a_wclk_p_r<27> a_wclk_p_r<28> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<58> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<58> A_BIST_DIN<58> A_BIST_EN a_blc_r<107> a_blc_r<106> a_blc_r<105> a_blc_r<104> a_blt_r<107> a_blt_r<106> a_blt_r<105> a_blt_r<104> A_BM<58> a_dclk_n_r<26> a_dclk_n_r<27> a_dclk_p_r<26> a_dclk_p_r<27> A_DOUT<58> A_DIN<58> a_rclk_n_r<26> a_rclk_n_r<27> a_rclk_p_r<26> a_rclk_p_r<27> a_tieh<58> a_wclk_n_r<26> a_wclk_n_r<27> a_wclk_p_r<26> a_wclk_p_r<27> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<57> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<57> A_BIST_DIN<57> A_BIST_EN a_blc_r<103> a_blc_r<102> a_blc_r<101> a_blc_r<100> a_blt_r<103> a_blt_r<102> a_blt_r<101> a_blt_r<100> A_BM<57> a_dclk_n_r<25> a_dclk_n_r<26> a_dclk_p_r<25> a_dclk_p_r<26> A_DOUT<57> A_DIN<57> a_rclk_n_r<25> a_rclk_n_r<26> a_rclk_p_r<25> a_rclk_p_r<26> a_tieh<57> a_wclk_n_r<25> a_wclk_n_r<26> a_wclk_p_r<25> a_wclk_p_r<26> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<56> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<56> A_BIST_DIN<56> A_BIST_EN a_blc_r<99> a_blc_r<98> a_blc_r<97> a_blc_r<96> a_blt_r<99> a_blt_r<98> a_blt_r<97> a_blt_r<96> A_BM<56> a_dclk_n_r<24> a_dclk_n_r<25> a_dclk_p_r<24> a_dclk_p_r<25> A_DOUT<56> A_DIN<56> a_rclk_n_r<24> a_rclk_n_r<25> a_rclk_p_r<24> a_rclk_p_r<25> a_tieh<56> a_wclk_n_r<24> a_wclk_n_r<25> a_wclk_p_r<24> a_wclk_p_r<25> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<55> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<55> A_BIST_DIN<55> A_BIST_EN a_blc_r<95> a_blc_r<94> a_blc_r<93> a_blc_r<92> a_blt_r<95> a_blt_r<94> a_blt_r<93> a_blt_r<92> A_BM<55> a_dclk_n_r<23> a_dclk_n_r<24> a_dclk_p_r<23> a_dclk_p_r<24> A_DOUT<55> A_DIN<55> a_rclk_n_r<23> a_rclk_n_r<24> a_rclk_p_r<23> a_rclk_p_r<24> a_tieh<55> a_wclk_n_r<23> a_wclk_n_r<24> a_wclk_p_r<23> a_wclk_p_r<24> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<54> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<54> A_BIST_DIN<54> A_BIST_EN a_blc_r<91> a_blc_r<90> a_blc_r<89> a_blc_r<88> a_blt_r<91> a_blt_r<90> a_blt_r<89> a_blt_r<88> A_BM<54> a_dclk_n_r<22> a_dclk_n_r<23> a_dclk_p_r<22> a_dclk_p_r<23> A_DOUT<54> A_DIN<54> a_rclk_n_r<22> a_rclk_n_r<23> a_rclk_p_r<22> a_rclk_p_r<23> a_tieh<54> a_wclk_n_r<22> a_wclk_n_r<23> a_wclk_p_r<22> a_wclk_p_r<23> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<53> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<53> A_BIST_DIN<53> A_BIST_EN a_blc_r<87> a_blc_r<86> a_blc_r<85> a_blc_r<84> a_blt_r<87> a_blt_r<86> a_blt_r<85> a_blt_r<84> A_BM<53> a_dclk_n_r<21> a_dclk_n_r<22> a_dclk_p_r<21> a_dclk_p_r<22> A_DOUT<53> A_DIN<53> a_rclk_n_r<21> a_rclk_n_r<22> a_rclk_p_r<21> a_rclk_p_r<22> a_tieh<53> a_wclk_n_r<21> a_wclk_n_r<22> a_wclk_p_r<21> a_wclk_p_r<22> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<52> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<52> A_BIST_DIN<52> A_BIST_EN a_blc_r<83> a_blc_r<82> a_blc_r<81> a_blc_r<80> a_blt_r<83> a_blt_r<82> a_blt_r<81> a_blt_r<80> A_BM<52> a_dclk_n_r<20> a_dclk_n_r<21> a_dclk_p_r<20> a_dclk_p_r<21> A_DOUT<52> A_DIN<52> a_rclk_n_r<20> a_rclk_n_r<21> a_rclk_p_r<20> a_rclk_p_r<21> a_tieh<52> a_wclk_n_r<20> a_wclk_n_r<21> a_wclk_p_r<20> a_wclk_p_r<21> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<51> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<51> A_BIST_DIN<51> A_BIST_EN a_blc_r<79> a_blc_r<78> a_blc_r<77> a_blc_r<76> a_blt_r<79> a_blt_r<78> a_blt_r<77> a_blt_r<76> A_BM<51> a_dclk_n_r<19> a_dclk_n_r<20> a_dclk_p_r<19> a_dclk_p_r<20> A_DOUT<51> A_DIN<51> a_rclk_n_r<19> a_rclk_n_r<20> a_rclk_p_r<19> a_rclk_p_r<20> a_tieh<51> a_wclk_n_r<19> a_wclk_n_r<20> a_wclk_p_r<19> a_wclk_p_r<20> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<50> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<50> A_BIST_DIN<50> A_BIST_EN a_blc_r<75> a_blc_r<74> a_blc_r<73> a_blc_r<72> a_blt_r<75> a_blt_r<74> a_blt_r<73> a_blt_r<72> A_BM<50> a_dclk_n_r<18> a_dclk_n_r<19> a_dclk_p_r<18> a_dclk_p_r<19> A_DOUT<50> A_DIN<50> a_rclk_n_r<18> a_rclk_n_r<19> a_rclk_p_r<18> a_rclk_p_r<19> a_tieh<50> a_wclk_n_r<18> a_wclk_n_r<19> a_wclk_p_r<18> a_wclk_p_r<19> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<49> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<49> A_BIST_DIN<49> A_BIST_EN a_blc_r<71> a_blc_r<70> a_blc_r<69> a_blc_r<68> a_blt_r<71> a_blt_r<70> a_blt_r<69> a_blt_r<68> A_BM<49> a_dclk_n_r<17> a_dclk_n_r<18> a_dclk_p_r<17> a_dclk_p_r<18> A_DOUT<49> A_DIN<49> a_rclk_n_r<17> a_rclk_n_r<18> a_rclk_p_r<17> a_rclk_p_r<18> a_tieh<49> a_wclk_n_r<17> a_wclk_n_r<18> a_wclk_p_r<17> a_wclk_p_r<18> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<48> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<48> A_BIST_DIN<48> A_BIST_EN a_blc_r<67> a_blc_r<66> a_blc_r<65> a_blc_r<64> a_blt_r<67> a_blt_r<66> a_blt_r<65> a_blt_r<64> A_BM<48> a_dclk_n_r<16> a_dclk_n_r<17> a_dclk_p_r<16> a_dclk_p_r<17> A_DOUT<48> A_DIN<48> a_rclk_n_r<16> a_rclk_n_r<17> a_rclk_p_r<16> a_rclk_p_r<17> a_tieh<48> a_wclk_n_r<16> a_wclk_n_r<17> a_wclk_p_r<16> a_wclk_p_r<17> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<47> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<47> A_BIST_DIN<47> A_BIST_EN a_blc_r<63> a_blc_r<62> a_blc_r<61> a_blc_r<60> a_blt_r<63> a_blt_r<62> a_blt_r<61> a_blt_r<60> A_BM<47> a_dclk_n_r<15> a_dclk_n_r<16> a_dclk_p_r<15> a_dclk_p_r<16> A_DOUT<47> A_DIN<47> a_rclk_n_r<15> a_rclk_n_r<16> a_rclk_p_r<15> a_rclk_p_r<16> a_tieh<47> a_wclk_n_r<15> a_wclk_n_r<16> a_wclk_p_r<15> a_wclk_p_r<16> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<46> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<46> A_BIST_DIN<46> A_BIST_EN a_blc_r<59> a_blc_r<58> a_blc_r<57> a_blc_r<56> a_blt_r<59> a_blt_r<58> a_blt_r<57> a_blt_r<56> A_BM<46> a_dclk_n_r<14> a_dclk_n_r<15> a_dclk_p_r<14> a_dclk_p_r<15> A_DOUT<46> A_DIN<46> a_rclk_n_r<14> a_rclk_n_r<15> a_rclk_p_r<14> a_rclk_p_r<15> a_tieh<46> a_wclk_n_r<14> a_wclk_n_r<15> a_wclk_p_r<14> a_wclk_p_r<15> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<45> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<45> A_BIST_DIN<45> A_BIST_EN a_blc_r<55> a_blc_r<54> a_blc_r<53> a_blc_r<52> a_blt_r<55> a_blt_r<54> a_blt_r<53> a_blt_r<52> A_BM<45> a_dclk_n_r<13> a_dclk_n_r<14> a_dclk_p_r<13> a_dclk_p_r<14> A_DOUT<45> A_DIN<45> a_rclk_n_r<13> a_rclk_n_r<14> a_rclk_p_r<13> a_rclk_p_r<14> a_tieh<45> a_wclk_n_r<13> a_wclk_n_r<14> a_wclk_p_r<13> a_wclk_p_r<14> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<44> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<44> A_BIST_DIN<44> A_BIST_EN a_blc_r<51> a_blc_r<50> a_blc_r<49> a_blc_r<48> a_blt_r<51> a_blt_r<50> a_blt_r<49> a_blt_r<48> A_BM<44> a_dclk_n_r<12> a_dclk_n_r<13> a_dclk_p_r<12> a_dclk_p_r<13> A_DOUT<44> A_DIN<44> a_rclk_n_r<12> a_rclk_n_r<13> a_rclk_p_r<12> a_rclk_p_r<13> a_tieh<44> a_wclk_n_r<12> a_wclk_n_r<13> a_wclk_p_r<12> a_wclk_p_r<13> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<43> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<43> A_BIST_DIN<43> A_BIST_EN a_blc_r<47> a_blc_r<46> a_blc_r<45> a_blc_r<44> a_blt_r<47> a_blt_r<46> a_blt_r<45> a_blt_r<44> A_BM<43> a_dclk_n_r<11> a_dclk_n_r<12> a_dclk_p_r<11> a_dclk_p_r<12> A_DOUT<43> A_DIN<43> a_rclk_n_r<11> a_rclk_n_r<12> a_rclk_p_r<11> a_rclk_p_r<12> a_tieh<43> a_wclk_n_r<11> a_wclk_n_r<12> a_wclk_p_r<11> a_wclk_p_r<12> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<42> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<42> A_BIST_DIN<42> A_BIST_EN a_blc_r<43> a_blc_r<42> a_blc_r<41> a_blc_r<40> a_blt_r<43> a_blt_r<42> a_blt_r<41> a_blt_r<40> A_BM<42> a_dclk_n_r<10> a_dclk_n_r<11> a_dclk_p_r<10> a_dclk_p_r<11> A_DOUT<42> A_DIN<42> a_rclk_n_r<10> a_rclk_n_r<11> a_rclk_p_r<10> a_rclk_p_r<11> a_tieh<42> a_wclk_n_r<10> a_wclk_n_r<11> a_wclk_p_r<10> a_wclk_p_r<11> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<41> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<41> A_BIST_DIN<41> A_BIST_EN a_blc_r<39> a_blc_r<38> a_blc_r<37> a_blc_r<36> a_blt_r<39> a_blt_r<38> a_blt_r<37> a_blt_r<36> A_BM<41> a_dclk_n_r<9> a_dclk_n_r<10> a_dclk_p_r<9> a_dclk_p_r<10> A_DOUT<41> A_DIN<41> a_rclk_n_r<9> a_rclk_n_r<10> a_rclk_p_r<9> a_rclk_p_r<10> a_tieh<41> a_wclk_n_r<9> a_wclk_n_r<10> a_wclk_p_r<9> a_wclk_p_r<10> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<40> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<40> A_BIST_DIN<40> A_BIST_EN a_blc_r<35> a_blc_r<34> a_blc_r<33> a_blc_r<32> a_blt_r<35> a_blt_r<34> a_blt_r<33> a_blt_r<32> A_BM<40> a_dclk_n_r<8> a_dclk_n_r<9> a_dclk_p_r<8> a_dclk_p_r<9> A_DOUT<40> A_DIN<40> a_rclk_n_r<8> a_rclk_n_r<9> a_rclk_p_r<8> a_rclk_p_r<9> a_tieh<40> a_wclk_n_r<8> a_wclk_n_r<9> a_wclk_p_r<8> a_wclk_p_r<9> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<39> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<39> A_BIST_DIN<39> A_BIST_EN a_blc_r<31> a_blc_r<30> a_blc_r<29> a_blc_r<28> a_blt_r<31> a_blt_r<30> a_blt_r<29> a_blt_r<28> A_BM<39> a_dclk_n_r<7> a_dclk_n_r<8> a_dclk_p_r<7> a_dclk_p_r<8> A_DOUT<39> A_DIN<39> a_rclk_n_r<7> a_rclk_n_r<8> a_rclk_p_r<7> a_rclk_p_r<8> a_tieh<39> a_wclk_n_r<7> a_wclk_n_r<8> a_wclk_p_r<7> a_wclk_p_r<8> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<38> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<38> A_BIST_DIN<38> A_BIST_EN a_blc_r<27> a_blc_r<26> a_blc_r<25> a_blc_r<24> a_blt_r<27> a_blt_r<26> a_blt_r<25> a_blt_r<24> A_BM<38> a_dclk_n_r<6> a_dclk_n_r<7> a_dclk_p_r<6> a_dclk_p_r<7> A_DOUT<38> A_DIN<38> a_rclk_n_r<6> a_rclk_n_r<7> a_rclk_p_r<6> a_rclk_p_r<7> a_tieh<38> a_wclk_n_r<6> a_wclk_n_r<7> a_wclk_p_r<6> a_wclk_p_r<7> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<37> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<37> A_BIST_DIN<37> A_BIST_EN a_blc_r<23> a_blc_r<22> a_blc_r<21> a_blc_r<20> a_blt_r<23> a_blt_r<22> a_blt_r<21> a_blt_r<20> A_BM<37> a_dclk_n_r<5> a_dclk_n_r<6> a_dclk_p_r<5> a_dclk_p_r<6> A_DOUT<37> A_DIN<37> a_rclk_n_r<5> a_rclk_n_r<6> a_rclk_p_r<5> a_rclk_p_r<6> a_tieh<37> a_wclk_n_r<5> a_wclk_n_r<6> a_wclk_p_r<5> a_wclk_p_r<6> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<36> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<36> A_BIST_DIN<36> A_BIST_EN a_blc_r<19> a_blc_r<18> a_blc_r<17> a_blc_r<16> a_blt_r<19> a_blt_r<18> a_blt_r<17> a_blt_r<16> A_BM<36> a_dclk_n_r<4> a_dclk_n_r<5> a_dclk_p_r<4> a_dclk_p_r<5> A_DOUT<36> A_DIN<36> a_rclk_n_r<4> a_rclk_n_r<5> a_rclk_p_r<4> a_rclk_p_r<5> a_tieh<36> a_wclk_n_r<4> a_wclk_n_r<5> a_wclk_p_r<4> a_wclk_p_r<5> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<35> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<35> A_BIST_DIN<35> A_BIST_EN a_blc_r<15> a_blc_r<14> a_blc_r<13> a_blc_r<12> a_blt_r<15> a_blt_r<14> a_blt_r<13> a_blt_r<12> A_BM<35> a_dclk_n_r<3> a_dclk_n_r<4> a_dclk_p_r<3> a_dclk_p_r<4> A_DOUT<35> A_DIN<35> a_rclk_n_r<3> a_rclk_n_r<4> a_rclk_p_r<3> a_rclk_p_r<4> a_tieh<35> a_wclk_n_r<3> a_wclk_n_r<4> a_wclk_p_r<3> a_wclk_p_r<4> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<34> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<34> A_BIST_DIN<34> A_BIST_EN a_blc_r<11> a_blc_r<10> a_blc_r<9> a_blc_r<8> a_blt_r<11> a_blt_r<10> a_blt_r<9> a_blt_r<8> A_BM<34> a_dclk_n_r<2> a_dclk_n_r<3> a_dclk_p_r<2> a_dclk_p_r<3> A_DOUT<34> A_DIN<34> a_rclk_n_r<2> a_rclk_n_r<3> a_rclk_p_r<2> a_rclk_p_r<3> a_tieh<34> a_wclk_n_r<2> a_wclk_n_r<3> a_wclk_p_r<2> a_wclk_p_r<3> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<33> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<33> A_BIST_DIN<33> A_BIST_EN a_blc_r<7> a_blc_r<6> a_blc_r<5> a_blc_r<4> a_blt_r<7> a_blt_r<6> a_blt_r<5> a_blt_r<4> A_BM<33> a_dclk_n_r<1> a_dclk_n_r<2> a_dclk_p_r<1> a_dclk_p_r<2> A_DOUT<33> A_DIN<33> a_rclk_n_r<1> a_rclk_n_r<2> a_rclk_p_r<1> a_rclk_p_r<2> a_tieh<33> a_wclk_n_r<1> a_wclk_n_r<2> a_wclk_p_r<1> a_wclk_p_r<2> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<32> a_addr_dec_r<3> a_addr_dec_r<2> a_addr_dec_r<1> a_addr_dec_r<0> A_BIST_BM<32> A_BIST_DIN<32> A_BIST_EN a_blc_r<3> a_blc_r<2> a_blc_r<1> a_blc_r<0> a_blt_r<3> a_blt_r<2> a_blt_r<1> a_blt_r<0> A_BM<32> a_dclk_n_r<0> a_dclk_n_r<1> a_dclk_p_r<0> a_dclk_p_r<1> A_DOUT<32> A_DIN<32> a_rclk_n_r<0> a_rclk_n_r<1> a_rclk_p_r<0> a_rclk_p_r<1> a_tieh<32> a_wclk_n_r<0> a_wclk_n_r<1> a_wclk_p_r<0> a_wclk_p_r<1> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<31> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<0> A_BIST_DIN<0> A_BIST_EN a_blc_l<127> a_blc_l<126> a_blc_l<125> a_blc_l<124> a_blt_l<127> a_blt_l<126> a_blt_l<125> a_blt_l<124> A_BM<0> a_dclk_n_l<31> a_dclk_n_l<32> a_dclk_p_l<31> a_dclk_p_l<32> A_DOUT<0> A_DIN<0> a_rclk_n_l<31> a_rclk_n_l<32> a_rclk_p_l<31> a_rclk_p_l<32> a_tieh<0> a_wclk_n_l<31> a_wclk_n_l<32> a_wclk_p_l<31> a_wclk_p_l<32> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<30> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<1> A_BIST_DIN<1> A_BIST_EN a_blc_l<123> a_blc_l<122> a_blc_l<121> a_blc_l<120> a_blt_l<123> a_blt_l<122> a_blt_l<121> a_blt_l<120> A_BM<1> a_dclk_n_l<30> a_dclk_n_l<31> a_dclk_p_l<30> a_dclk_p_l<31> A_DOUT<1> A_DIN<1> a_rclk_n_l<30> a_rclk_n_l<31> a_rclk_p_l<30> a_rclk_p_l<31> a_tieh<1> a_wclk_n_l<30> a_wclk_n_l<31> a_wclk_p_l<30> a_wclk_p_l<31> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<29> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<2> A_BIST_DIN<2> A_BIST_EN a_blc_l<119> a_blc_l<118> a_blc_l<117> a_blc_l<116> a_blt_l<119> a_blt_l<118> a_blt_l<117> a_blt_l<116> A_BM<2> a_dclk_n_l<29> a_dclk_n_l<30> a_dclk_p_l<29> a_dclk_p_l<30> A_DOUT<2> A_DIN<2> a_rclk_n_l<29> a_rclk_n_l<30> a_rclk_p_l<29> a_rclk_p_l<30> a_tieh<2> a_wclk_n_l<29> a_wclk_n_l<30> a_wclk_p_l<29> a_wclk_p_l<30> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<28> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<3> A_BIST_DIN<3> A_BIST_EN a_blc_l<115> a_blc_l<114> a_blc_l<113> a_blc_l<112> a_blt_l<115> a_blt_l<114> a_blt_l<113> a_blt_l<112> A_BM<3> a_dclk_n_l<28> a_dclk_n_l<29> a_dclk_p_l<28> a_dclk_p_l<29> A_DOUT<3> A_DIN<3> a_rclk_n_l<28> a_rclk_n_l<29> a_rclk_p_l<28> a_rclk_p_l<29> a_tieh<3> a_wclk_n_l<28> a_wclk_n_l<29> a_wclk_p_l<28> a_wclk_p_l<29> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<27> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<4> A_BIST_DIN<4> A_BIST_EN a_blc_l<111> a_blc_l<110> a_blc_l<109> a_blc_l<108> a_blt_l<111> a_blt_l<110> a_blt_l<109> a_blt_l<108> A_BM<4> a_dclk_n_l<27> a_dclk_n_l<28> a_dclk_p_l<27> a_dclk_p_l<28> A_DOUT<4> A_DIN<4> a_rclk_n_l<27> a_rclk_n_l<28> a_rclk_p_l<27> a_rclk_p_l<28> a_tieh<4> a_wclk_n_l<27> a_wclk_n_l<28> a_wclk_p_l<27> a_wclk_p_l<28> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<26> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<5> A_BIST_DIN<5> A_BIST_EN a_blc_l<107> a_blc_l<106> a_blc_l<105> a_blc_l<104> a_blt_l<107> a_blt_l<106> a_blt_l<105> a_blt_l<104> A_BM<5> a_dclk_n_l<26> a_dclk_n_l<27> a_dclk_p_l<26> a_dclk_p_l<27> A_DOUT<5> A_DIN<5> a_rclk_n_l<26> a_rclk_n_l<27> a_rclk_p_l<26> a_rclk_p_l<27> a_tieh<5> a_wclk_n_l<26> a_wclk_n_l<27> a_wclk_p_l<26> a_wclk_p_l<27> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<25> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<6> A_BIST_DIN<6> A_BIST_EN a_blc_l<103> a_blc_l<102> a_blc_l<101> a_blc_l<100> a_blt_l<103> a_blt_l<102> a_blt_l<101> a_blt_l<100> A_BM<6> a_dclk_n_l<25> a_dclk_n_l<26> a_dclk_p_l<25> a_dclk_p_l<26> A_DOUT<6> A_DIN<6> a_rclk_n_l<25> a_rclk_n_l<26> a_rclk_p_l<25> a_rclk_p_l<26> a_tieh<6> a_wclk_n_l<25> a_wclk_n_l<26> a_wclk_p_l<25> a_wclk_p_l<26> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<24> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<7> A_BIST_DIN<7> A_BIST_EN a_blc_l<99> a_blc_l<98> a_blc_l<97> a_blc_l<96> a_blt_l<99> a_blt_l<98> a_blt_l<97> a_blt_l<96> A_BM<7> a_dclk_n_l<24> a_dclk_n_l<25> a_dclk_p_l<24> a_dclk_p_l<25> A_DOUT<7> A_DIN<7> a_rclk_n_l<24> a_rclk_n_l<25> a_rclk_p_l<24> a_rclk_p_l<25> a_tieh<7> a_wclk_n_l<24> a_wclk_n_l<25> a_wclk_p_l<24> a_wclk_p_l<25> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<23> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<8> A_BIST_DIN<8> A_BIST_EN a_blc_l<95> a_blc_l<94> a_blc_l<93> a_blc_l<92> a_blt_l<95> a_blt_l<94> a_blt_l<93> a_blt_l<92> A_BM<8> a_dclk_n_l<23> a_dclk_n_l<24> a_dclk_p_l<23> a_dclk_p_l<24> A_DOUT<8> A_DIN<8> a_rclk_n_l<23> a_rclk_n_l<24> a_rclk_p_l<23> a_rclk_p_l<24> a_tieh<8> a_wclk_n_l<23> a_wclk_n_l<24> a_wclk_p_l<23> a_wclk_p_l<24> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<22> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<9> A_BIST_DIN<9> A_BIST_EN a_blc_l<91> a_blc_l<90> a_blc_l<89> a_blc_l<88> a_blt_l<91> a_blt_l<90> a_blt_l<89> a_blt_l<88> A_BM<9> a_dclk_n_l<22> a_dclk_n_l<23> a_dclk_p_l<22> a_dclk_p_l<23> A_DOUT<9> A_DIN<9> a_rclk_n_l<22> a_rclk_n_l<23> a_rclk_p_l<22> a_rclk_p_l<23> a_tieh<9> a_wclk_n_l<22> a_wclk_n_l<23> a_wclk_p_l<22> a_wclk_p_l<23> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<21> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<10> A_BIST_DIN<10> A_BIST_EN a_blc_l<87> a_blc_l<86> a_blc_l<85> a_blc_l<84> a_blt_l<87> a_blt_l<86> a_blt_l<85> a_blt_l<84> A_BM<10> a_dclk_n_l<21> a_dclk_n_l<22> a_dclk_p_l<21> a_dclk_p_l<22> A_DOUT<10> A_DIN<10> a_rclk_n_l<21> a_rclk_n_l<22> a_rclk_p_l<21> a_rclk_p_l<22> a_tieh<10> a_wclk_n_l<21> a_wclk_n_l<22> a_wclk_p_l<21> a_wclk_p_l<22> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<20> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<11> A_BIST_DIN<11> A_BIST_EN a_blc_l<83> a_blc_l<82> a_blc_l<81> a_blc_l<80> a_blt_l<83> a_blt_l<82> a_blt_l<81> a_blt_l<80> A_BM<11> a_dclk_n_l<20> a_dclk_n_l<21> a_dclk_p_l<20> a_dclk_p_l<21> A_DOUT<11> A_DIN<11> a_rclk_n_l<20> a_rclk_n_l<21> a_rclk_p_l<20> a_rclk_p_l<21> a_tieh<11> a_wclk_n_l<20> a_wclk_n_l<21> a_wclk_p_l<20> a_wclk_p_l<21> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<19> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<12> A_BIST_DIN<12> A_BIST_EN a_blc_l<79> a_blc_l<78> a_blc_l<77> a_blc_l<76> a_blt_l<79> a_blt_l<78> a_blt_l<77> a_blt_l<76> A_BM<12> a_dclk_n_l<19> a_dclk_n_l<20> a_dclk_p_l<19> a_dclk_p_l<20> A_DOUT<12> A_DIN<12> a_rclk_n_l<19> a_rclk_n_l<20> a_rclk_p_l<19> a_rclk_p_l<20> a_tieh<12> a_wclk_n_l<19> a_wclk_n_l<20> a_wclk_p_l<19> a_wclk_p_l<20> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<18> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<13> A_BIST_DIN<13> A_BIST_EN a_blc_l<75> a_blc_l<74> a_blc_l<73> a_blc_l<72> a_blt_l<75> a_blt_l<74> a_blt_l<73> a_blt_l<72> A_BM<13> a_dclk_n_l<18> a_dclk_n_l<19> a_dclk_p_l<18> a_dclk_p_l<19> A_DOUT<13> A_DIN<13> a_rclk_n_l<18> a_rclk_n_l<19> a_rclk_p_l<18> a_rclk_p_l<19> a_tieh<13> a_wclk_n_l<18> a_wclk_n_l<19> a_wclk_p_l<18> a_wclk_p_l<19> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<17> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<14> A_BIST_DIN<14> A_BIST_EN a_blc_l<71> a_blc_l<70> a_blc_l<69> a_blc_l<68> a_blt_l<71> a_blt_l<70> a_blt_l<69> a_blt_l<68> A_BM<14> a_dclk_n_l<17> a_dclk_n_l<18> a_dclk_p_l<17> a_dclk_p_l<18> A_DOUT<14> A_DIN<14> a_rclk_n_l<17> a_rclk_n_l<18> a_rclk_p_l<17> a_rclk_p_l<18> a_tieh<14> a_wclk_n_l<17> a_wclk_n_l<18> a_wclk_p_l<17> a_wclk_p_l<18> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<16> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<15> A_BIST_DIN<15> A_BIST_EN a_blc_l<67> a_blc_l<66> a_blc_l<65> a_blc_l<64> a_blt_l<67> a_blt_l<66> a_blt_l<65> a_blt_l<64> A_BM<15> a_dclk_n_l<16> a_dclk_n_l<17> a_dclk_p_l<16> a_dclk_p_l<17> A_DOUT<15> A_DIN<15> a_rclk_n_l<16> a_rclk_n_l<17> a_rclk_p_l<16> a_rclk_p_l<17> a_tieh<15> a_wclk_n_l<16> a_wclk_n_l<17> a_wclk_p_l<16> a_wclk_p_l<17> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<15> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<16> A_BIST_DIN<16> A_BIST_EN a_blc_l<63> a_blc_l<62> a_blc_l<61> a_blc_l<60> a_blt_l<63> a_blt_l<62> a_blt_l<61> a_blt_l<60> A_BM<16> a_dclk_n_l<15> a_dclk_n_l<16> a_dclk_p_l<15> a_dclk_p_l<16> A_DOUT<16> A_DIN<16> a_rclk_n_l<15> a_rclk_n_l<16> a_rclk_p_l<15> a_rclk_p_l<16> a_tieh<16> a_wclk_n_l<15> a_wclk_n_l<16> a_wclk_p_l<15> a_wclk_p_l<16> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<14> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<17> A_BIST_DIN<17> A_BIST_EN a_blc_l<59> a_blc_l<58> a_blc_l<57> a_blc_l<56> a_blt_l<59> a_blt_l<58> a_blt_l<57> a_blt_l<56> A_BM<17> a_dclk_n_l<14> a_dclk_n_l<15> a_dclk_p_l<14> a_dclk_p_l<15> A_DOUT<17> A_DIN<17> a_rclk_n_l<14> a_rclk_n_l<15> a_rclk_p_l<14> a_rclk_p_l<15> a_tieh<17> a_wclk_n_l<14> a_wclk_n_l<15> a_wclk_p_l<14> a_wclk_p_l<15> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<13> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<18> A_BIST_DIN<18> A_BIST_EN a_blc_l<55> a_blc_l<54> a_blc_l<53> a_blc_l<52> a_blt_l<55> a_blt_l<54> a_blt_l<53> a_blt_l<52> A_BM<18> a_dclk_n_l<13> a_dclk_n_l<14> a_dclk_p_l<13> a_dclk_p_l<14> A_DOUT<18> A_DIN<18> a_rclk_n_l<13> a_rclk_n_l<14> a_rclk_p_l<13> a_rclk_p_l<14> a_tieh<18> a_wclk_n_l<13> a_wclk_n_l<14> a_wclk_p_l<13> a_wclk_p_l<14> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<12> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<19> A_BIST_DIN<19> A_BIST_EN a_blc_l<51> a_blc_l<50> a_blc_l<49> a_blc_l<48> a_blt_l<51> a_blt_l<50> a_blt_l<49> a_blt_l<48> A_BM<19> a_dclk_n_l<12> a_dclk_n_l<13> a_dclk_p_l<12> a_dclk_p_l<13> A_DOUT<19> A_DIN<19> a_rclk_n_l<12> a_rclk_n_l<13> a_rclk_p_l<12> a_rclk_p_l<13> a_tieh<19> a_wclk_n_l<12> a_wclk_n_l<13> a_wclk_p_l<12> a_wclk_p_l<13> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<11> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<20> A_BIST_DIN<20> A_BIST_EN a_blc_l<47> a_blc_l<46> a_blc_l<45> a_blc_l<44> a_blt_l<47> a_blt_l<46> a_blt_l<45> a_blt_l<44> A_BM<20> a_dclk_n_l<11> a_dclk_n_l<12> a_dclk_p_l<11> a_dclk_p_l<12> A_DOUT<20> A_DIN<20> a_rclk_n_l<11> a_rclk_n_l<12> a_rclk_p_l<11> a_rclk_p_l<12> a_tieh<20> a_wclk_n_l<11> a_wclk_n_l<12> a_wclk_p_l<11> a_wclk_p_l<12> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<10> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<21> A_BIST_DIN<21> A_BIST_EN a_blc_l<43> a_blc_l<42> a_blc_l<41> a_blc_l<40> a_blt_l<43> a_blt_l<42> a_blt_l<41> a_blt_l<40> A_BM<21> a_dclk_n_l<10> a_dclk_n_l<11> a_dclk_p_l<10> a_dclk_p_l<11> A_DOUT<21> A_DIN<21> a_rclk_n_l<10> a_rclk_n_l<11> a_rclk_p_l<10> a_rclk_p_l<11> a_tieh<21> a_wclk_n_l<10> a_wclk_n_l<11> a_wclk_p_l<10> a_wclk_p_l<11> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<9> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<22> A_BIST_DIN<22> A_BIST_EN a_blc_l<39> a_blc_l<38> a_blc_l<37> a_blc_l<36> a_blt_l<39> a_blt_l<38> a_blt_l<37> a_blt_l<36> A_BM<22> a_dclk_n_l<9> a_dclk_n_l<10> a_dclk_p_l<9> a_dclk_p_l<10> A_DOUT<22> A_DIN<22> a_rclk_n_l<9> a_rclk_n_l<10> a_rclk_p_l<9> a_rclk_p_l<10> a_tieh<22> a_wclk_n_l<9> a_wclk_n_l<10> a_wclk_p_l<9> a_wclk_p_l<10> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<8> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<23> A_BIST_DIN<23> A_BIST_EN a_blc_l<35> a_blc_l<34> a_blc_l<33> a_blc_l<32> a_blt_l<35> a_blt_l<34> a_blt_l<33> a_blt_l<32> A_BM<23> a_dclk_n_l<8> a_dclk_n_l<9> a_dclk_p_l<8> a_dclk_p_l<9> A_DOUT<23> A_DIN<23> a_rclk_n_l<8> a_rclk_n_l<9> a_rclk_p_l<8> a_rclk_p_l<9> a_tieh<23> a_wclk_n_l<8> a_wclk_n_l<9> a_wclk_p_l<8> a_wclk_p_l<9> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<7> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<24> A_BIST_DIN<24> A_BIST_EN a_blc_l<31> a_blc_l<30> a_blc_l<29> a_blc_l<28> a_blt_l<31> a_blt_l<30> a_blt_l<29> a_blt_l<28> A_BM<24> a_dclk_n_l<7> a_dclk_n_l<8> a_dclk_p_l<7> a_dclk_p_l<8> A_DOUT<24> A_DIN<24> a_rclk_n_l<7> a_rclk_n_l<8> a_rclk_p_l<7> a_rclk_p_l<8> a_tieh<24> a_wclk_n_l<7> a_wclk_n_l<8> a_wclk_p_l<7> a_wclk_p_l<8> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<6> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<25> A_BIST_DIN<25> A_BIST_EN a_blc_l<27> a_blc_l<26> a_blc_l<25> a_blc_l<24> a_blt_l<27> a_blt_l<26> a_blt_l<25> a_blt_l<24> A_BM<25> a_dclk_n_l<6> a_dclk_n_l<7> a_dclk_p_l<6> a_dclk_p_l<7> A_DOUT<25> A_DIN<25> a_rclk_n_l<6> a_rclk_n_l<7> a_rclk_p_l<6> a_rclk_p_l<7> a_tieh<25> a_wclk_n_l<6> a_wclk_n_l<7> a_wclk_p_l<6> a_wclk_p_l<7> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<5> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<26> A_BIST_DIN<26> A_BIST_EN a_blc_l<23> a_blc_l<22> a_blc_l<21> a_blc_l<20> a_blt_l<23> a_blt_l<22> a_blt_l<21> a_blt_l<20> A_BM<26> a_dclk_n_l<5> a_dclk_n_l<6> a_dclk_p_l<5> a_dclk_p_l<6> A_DOUT<26> A_DIN<26> a_rclk_n_l<5> a_rclk_n_l<6> a_rclk_p_l<5> a_rclk_p_l<6> a_tieh<26> a_wclk_n_l<5> a_wclk_n_l<6> a_wclk_p_l<5> a_wclk_p_l<6> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<4> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<27> A_BIST_DIN<27> A_BIST_EN a_blc_l<19> a_blc_l<18> a_blc_l<17> a_blc_l<16> a_blt_l<19> a_blt_l<18> a_blt_l<17> a_blt_l<16> A_BM<27> a_dclk_n_l<4> a_dclk_n_l<5> a_dclk_p_l<4> a_dclk_p_l<5> A_DOUT<27> A_DIN<27> a_rclk_n_l<4> a_rclk_n_l<5> a_rclk_p_l<4> a_rclk_p_l<5> a_tieh<27> a_wclk_n_l<4> a_wclk_n_l<5> a_wclk_p_l<4> a_wclk_p_l<5> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<3> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<28> A_BIST_DIN<28> A_BIST_EN a_blc_l<15> a_blc_l<14> a_blc_l<13> a_blc_l<12> a_blt_l<15> a_blt_l<14> a_blt_l<13> a_blt_l<12> A_BM<28> a_dclk_n_l<3> a_dclk_n_l<4> a_dclk_p_l<3> a_dclk_p_l<4> A_DOUT<28> A_DIN<28> a_rclk_n_l<3> a_rclk_n_l<4> a_rclk_p_l<3> a_rclk_p_l<4> a_tieh<28> a_wclk_n_l<3> a_wclk_n_l<4> a_wclk_p_l<3> a_wclk_p_l<4> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<2> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<29> A_BIST_DIN<29> A_BIST_EN a_blc_l<11> a_blc_l<10> a_blc_l<9> a_blc_l<8> a_blt_l<11> a_blt_l<10> a_blt_l<9> a_blt_l<8> A_BM<29> a_dclk_n_l<2> a_dclk_n_l<3> a_dclk_p_l<2> a_dclk_p_l<3> A_DOUT<29> A_DIN<29> a_rclk_n_l<2> a_rclk_n_l<3> a_rclk_p_l<2> a_rclk_p_l<3> a_tieh<29> a_wclk_n_l<2> a_wclk_n_l<3> a_wclk_p_l<2> a_wclk_p_l<3> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<1> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<30> A_BIST_DIN<30> A_BIST_EN a_blc_l<7> a_blc_l<6> a_blc_l<5> a_blc_l<4> a_blt_l<7> a_blt_l<6> a_blt_l<5> a_blt_l<4> A_BM<30> a_dclk_n_l<1> a_dclk_n_l<2> a_dclk_p_l<1> a_dclk_p_l<2> A_DOUT<30> A_DIN<30> a_rclk_n_l<1> a_rclk_n_l<2> a_rclk_p_l<1> a_rclk_p_l<2> a_tieh<30> a_wclk_n_l<1> a_wclk_n_l<2> a_wclk_p_l<1> a_wclk_p_l<2> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2
XCOLCTRL<0> a_addr_dec_l<3> a_addr_dec_l<2> a_addr_dec_l<1> a_addr_dec_l<0> A_BIST_BM<31> A_BIST_DIN<31> A_BIST_EN a_blc_l<3> a_blc_l<2> a_blc_l<1> a_blc_l<0> a_blt_l<3> a_blt_l<2> a_blt_l<1> a_blt_l<0> A_BM<31> a_dclk_n_l<0> a_dclk_n_l<1> a_dclk_p_l<0> a_dclk_p_l<1> A_DOUT<31> A_DIN<31> a_rclk_n_l<0> a_rclk_n_l<1> a_rclk_p_l<0> a_rclk_p_l<1> a_tieh<31> a_wclk_n_l<0> a_wclk_n_l<1> a_wclk_p_l<0> a_wclk_p_l<1> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLCTRL2


XDRVFILL4<1> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4
XDRVFILL4<2> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4
XDRVFILL4<3> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4
XDRVFILL4<4> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4
XCOLFILL4<1> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<2> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<3> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<4> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<5> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<6> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<7> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<8> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<9> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
XCOLFILL4<10> VDD! VSS! / RM_IHPSG13_2048x64_c2_1P_COLDRV13_FILL4C2
.ENDS
