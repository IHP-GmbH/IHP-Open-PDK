*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT inductor
L1 net1 net2 sub inductor w=2u s=2.1u d=25.35u nr_r=1
L2 net3 net4 sub inductor w=2u s=2.1u d=25.35u nr_r=2
L4 net5 net6 sub inductor w=2u s=2.1u d=25.35u nr_r=1
L5 net6 net5 sub inductor w=2u s=2.1u d=25.35u nr_r=1

* Extra patterns
L_pattern_1  la_1  lb_1  sub inductor w=8.22u s=3.29u d=47.65u nr_r=1 
L_pattern_2  la_2  lb_2  sub inductor w=9.34u s=3.29u d=53.06u nr_r=1 
L_pattern_3  la_3  lb_3  sub inductor w=5.42u s=5.73u d=40.02u nr_r=1 
L_pattern_4  la_4  lb_4  sub inductor w=5.34u s=8.97u d=47.45u nr_r=1 
L_pattern_5  la_5  lb_5  sub inductor w=5.42u s=3.74u d=48.39u nr_r=1 
L_pattern_6  la_6  lb_6  sub inductor w=7.0u s=3.74u d=45.33u nr_r=1 
L_pattern_7  la_7  lb_7  sub inductor w=3.31u s=4.29u d=25.63u nr_r=1 
L_pattern_8  la_8  lb_8  sub inductor w=6.1u s=7.11u d=48.39u nr_r=1 
L_pattern_9  la_9  lb_9  sub inductor w=2.6u s=4.29u d=33.29u nr_r=1 
L_pattern_10 la_10 lb_10 sub inductor w=2.6u s=3.73u d=25.63u nr_r=1 
L_pattern_11 la_11 lb_11 sub inductor w=8.22u s=3.74u d=141.975u nr_r=4
L_pattern_12 la_12 lb_12 sub inductor w=9.34u s=3.74u d=156.61u nr_r=4 
L_pattern_13 la_13 lb_13 sub inductor w=6.1u s=3.29u d=110.11u nr_r=5
L_pattern_14 la_14 lb_14 sub inductor w=5.42u s=4.29u d=110.47u nr_r=5 
L_pattern_15 la_15 lb_15 sub inductor w=5.34u s=5.73u d=122.735u nr_r=3
L_pattern_16 la_16 lb_16 sub inductor w=5.42u s=8.97u d=153.735u nr_r=3   
.ENDS
