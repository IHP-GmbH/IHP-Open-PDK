VBIC Gummel Test Ic=f(Vc,Vb)

.lib ../models/cornerHBT.lib hbt_typ

vb b 0 0.5
vc c 0 1.0
vs s 0 0.0
XQ1 C B 0 S t npn13G2 nx=1

.dc vb 0.2 1.2 0.01
.print dc v(b) i(vc) i(vb) i(vs)

.end
