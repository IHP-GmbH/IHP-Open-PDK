*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT dpantenna
D1 net1 VDD dpantenna w=780.00n l=780.00n a=608.400f p=3.12u m=1
D2 net2 VDD dpantenna w=800.00n l=780.00n a=624.000f p=3.16u m=1
D3 net3 VDD dpantenna w=780.00n l=700.00n a=546.000f p=2.96u m=1
D4 net4 VDD dpantenna w=780.00n l=780.00n a=608.400f p=3.12u m=2

* Extra patterns
D_pattern_1  anode_1  WELL dpantenna w=3.42u l=9.15u 
D_pattern_2  anode_2  WELL dpantenna w=2.91u l=8.9u 
D_pattern_3  anode_3  WELL dpantenna w=1.45u l=1.38u 
D_pattern_4  anode_4  WELL dpantenna w=2.03u l=7.77u 
D_pattern_5  anode_5  WELL dpantenna w=2.05u l=8.12u 
D_pattern_6  anode_6  WELL dpantenna w=3.87u l=4.67u 
D_pattern_7  anode_7  WELL dpantenna w=6.24u l=1.21u 
D_pattern_8  anode_8  WELL dpantenna w=9.78u l=6.53u 
D_pattern_9  anode_9  WELL dpantenna w=9.78u l=1.21u 
D_pattern_10 anode_10 WELL dpantenna w=6.24u l=4.67u 
D_pattern_11 anode_11 WELL dpantenna w=3.87u l=8.12u 
D_pattern_12 anode_12 WELL dpantenna w=2.05u l=7.77u 
D_pattern_13 anode_13 WELL dpantenna w=2.03u l=1.38u 
D_pattern_14 anode_14 WELL dpantenna w=1.45u l=8.9u 
D_pattern_15 anode_15 WELL dpantenna w=2.91u l=9.15u 
D_pattern_16 anode_16 WELL dpantenna w=3.42u l=6.53u 
D_pattern_17 anode_17 WELL dpantenna w=3.42u l=1.21u 
D_pattern_18 anode_18 WELL dpantenna w=2.91u l=4.67u 
D_pattern_19 anode_19 WELL dpantenna w=1.45u l=8.12u 
D_pattern_20 anode_20 WELL dpantenna w=2.03u l=6.53u 
D_pattern_21 anode_21 WELL dpantenna w=2.05u l=9.15u 
D_pattern_22 anode_22 WELL dpantenna w=3.87u l=8.9u 
D_pattern_23 anode_23 WELL dpantenna w=6.24u l=1.38u 
D_pattern_24 anode_24 WELL dpantenna w=9.78u l=7.77u 
D_pattern_25 anode_25 WELL dpantenna w=9.78u l=1.38u 
D_pattern_26 anode_26 WELL dpantenna w=6.24u l=8.9u 
D_pattern_27 anode_27 WELL dpantenna w=3.87u l=9.15u 
D_pattern_28 anode_28 WELL dpantenna w=2.05u l=6.53u 
D_pattern_29 anode_29 WELL dpantenna w=2.03u l=1.21u 
D_pattern_30 anode_30 WELL dpantenna w=1.45u l=4.67u 
D_pattern_31 anode_31 WELL dpantenna w=2.91u l=7.77u 
D_pattern_32 anode_32 WELL dpantenna w=3.42u l=8.12u 
D_pattern_33 anode_33 WELL dpantenna w=3.42u l=7.77u 
D_pattern_34 anode_34 WELL dpantenna w=2.91u l=1.38u 
D_pattern_35 anode_35 WELL dpantenna w=1.45u l=1.21u 
D_pattern_36 anode_36 WELL dpantenna w=2.03u l=9.15u 
D_pattern_37 anode_37 WELL dpantenna w=2.05u l=4.67u 
D_pattern_38 anode_38 WELL dpantenna w=3.87u l=6.53u 
D_pattern_39 anode_39 WELL dpantenna w=6.24u l=8.12u 
D_pattern_40 anode_40 WELL dpantenna w=9.78u l=8.9u 
D_pattern_41 anode_41 WELL dpantenna w=9.78u l=8.12u 
D_pattern_42 anode_42 WELL dpantenna w=6.24u l=9.15u 
D_pattern_43 anode_43 WELL dpantenna w=3.87u l=7.77u 
D_pattern_44 anode_44 WELL dpantenna w=2.05u l=1.21u 
D_pattern_45 anode_45 WELL dpantenna w=2.03u l=8.9u 
D_pattern_46 anode_46 WELL dpantenna w=1.45u l=6.53u 
D_pattern_47 anode_47 WELL dpantenna w=2.91u l=6.53u 
D_pattern_48 anode_48 WELL dpantenna w=3.42u l=4.67u 
D_pattern_49 anode_49 WELL dpantenna w=3.42u l=1.38u 
D_pattern_50 anode_50 WELL dpantenna w=2.91u l=8.12u 
D_pattern_51 anode_51 WELL dpantenna w=1.45u l=7.77u 
D_pattern_52 anode_52 WELL dpantenna w=2.03u l=4.67u 
D_pattern_53 anode_53 WELL dpantenna w=2.05u l=1.38u 
D_pattern_54 anode_54 WELL dpantenna w=3.87u l=1.21u 
D_pattern_55 anode_55 WELL dpantenna w=6.24u l=7.77u 
D_pattern_56 anode_56 WELL dpantenna w=9.78u l=9.15u 
D_pattern_57 anode_57 WELL dpantenna w=9.78u l=4.67u 
D_pattern_58 anode_58 WELL dpantenna w=6.24u l=6.53u 
D_pattern_59 anode_59 WELL dpantenna w=3.87u l=1.38u 
D_pattern_60 anode_60 WELL dpantenna w=2.05u l=8.9u 
D_pattern_61 anode_61 WELL dpantenna w=2.03u l=8.12u 
D_pattern_62 anode_62 WELL dpantenna w=1.45u l=9.15u 
D_pattern_63 anode_63 WELL dpantenna w=2.91u l=1.21u 
D_pattern_64 anode_64 WELL dpantenna w=3.42u l=8.9u 
D_pattern_65 anode_65 WELL dpantenna w=2.03u l=1.21u 
D_pattern_66 anode_66 WELL dpantenna w=3.87u l=6.53u 
.ENDS
