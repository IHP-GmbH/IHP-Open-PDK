psp103 test circuit
*
vd  d 0 dc 0.1
vg  g 0 dc 0.0
vs  s 0 dc 0.0
vb  b 0 dc 0.0
X1  d g s b sg13_lv_nmos w=1u l=0.13u mult=1
.option temp=21
.step  vb -3 0 0.5
.dc vg 0 1.5 0.02
.print dc format=gnuplot v(g) i(vd)
*
.lib ../models/cornerMOSlv.lib mos_tt

.end

