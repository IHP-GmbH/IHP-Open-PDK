*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT ntap1
R1 net1 WELL1 ntap1 A=608.4f Perim=3.12u
R2 net2 WELL2  ntap1 A=624.0f P=3.16u
R3 net3 WELL2  ntap1 A=640.0f P=3.20u

* Extra patterns
R_pattern_1  a_1  WELL ntap1 w=8.06u l=8.97u 
R_pattern_2  a_2  WELL ntap1 w=9.79u l=8.97u 
R_pattern_3  a_3  WELL ntap1 w=5.31u l=8.97u 
R_pattern_4  a_4  WELL ntap1 w=6.88u l=8.97u 
R_pattern_5  a_5  WELL ntap1 w=4.25u l=8.97u 
R_pattern_6  a_6  WELL ntap1 w=3.76u l=8.97u 
R_pattern_7  a_7  WELL ntap1 w=3.61u l=8.97u 
R_pattern_8  a_8  WELL ntap1 w=6.43u l=8.97u 
R_pattern_9  a_9  WELL ntap1 w=6.43u l=2.43u 
R_pattern_10 a_10 WELL ntap1 w=3.61u l=2.43u 
R_pattern_11 a_11 WELL ntap1 w=3.76u l=2.43u 
R_pattern_12 a_12 WELL ntap1 w=4.25u l=2.43u 
R_pattern_13 a_13 WELL ntap1 w=6.88u l=2.43u 
R_pattern_14 a_14 WELL ntap1 w=5.31u l=2.43u 
R_pattern_15 a_15 WELL ntap1 w=9.79u l=2.43u 
R_pattern_16 a_16 WELL ntap1 w=8.06u l=2.43u 
R_pattern_17 a_17 WELL ntap1 w=8.06u l=5.71u 
R_pattern_18 a_18 WELL ntap1 w=9.79u l=5.71u 
R_pattern_19 a_19 WELL ntap1 w=5.31u l=5.71u 
R_pattern_20 a_20 WELL ntap1 w=6.88u l=5.71u 
R_pattern_21 a_21 WELL ntap1 w=4.25u l=5.71u 
R_pattern_22 a_22 WELL ntap1 w=3.76u l=5.71u 
R_pattern_23 a_23 WELL ntap1 w=3.61u l=5.71u 
R_pattern_24 a_24 WELL ntap1 w=6.43u l=5.71u 
R_pattern_25 a_25 WELL ntap1 w=6.43u l=3.21u 
R_pattern_26 a_26 WELL ntap1 w=3.61u l=3.21u 
R_pattern_27 a_27 WELL ntap1 w=3.76u l=3.21u 
R_pattern_28 a_28 WELL ntap1 w=4.25u l=3.21u 
R_pattern_29 a_29 WELL ntap1 w=6.88u l=3.21u 
R_pattern_30 a_30 WELL ntap1 w=5.31u l=3.21u 
R_pattern_31 a_31 WELL ntap1 w=9.79u l=3.21u 
R_pattern_32 a_32 WELL ntap1 w=8.06u l=3.21u 
R_pattern_33 a_33 WELL ntap1 w=8.06u l=3.99u 
R_pattern_34 a_34 WELL ntap1 w=9.79u l=3.99u 
R_pattern_35 a_35 WELL ntap1 w=5.31u l=3.99u 
R_pattern_36 a_36 WELL ntap1 w=6.88u l=3.99u 
R_pattern_37 a_37 WELL ntap1 w=4.25u l=3.99u 
R_pattern_38 a_38 WELL ntap1 w=3.76u l=3.99u 
R_pattern_39 a_39 WELL ntap1 w=3.61u l=3.99u 
R_pattern_40 a_40 WELL ntap1 w=6.43u l=3.99u 
R_pattern_41 a_41 WELL ntap1 w=6.43u l=0.79u 
R_pattern_42 a_42 WELL ntap1 w=3.61u l=0.79u 
R_pattern_43 a_43 WELL ntap1 w=3.76u l=0.79u 
R_pattern_44 a_44 WELL ntap1 w=4.25u l=0.79u 
R_pattern_45 a_45 WELL ntap1 w=6.88u l=0.79u 
R_pattern_46 a_46 WELL ntap1 w=5.31u l=0.79u 
R_pattern_47 a_47 WELL ntap1 w=9.79u l=0.79u 
R_pattern_48 a_48 WELL ntap1 w=8.06u l=0.79u 
R_pattern_49 a_49 WELL ntap1 w=8.06u l=6.28u 
R_pattern_50 a_50 WELL ntap1 w=9.79u l=6.28u 
R_pattern_51 a_51 WELL ntap1 w=5.31u l=6.28u 
R_pattern_52 a_52 WELL ntap1 w=6.88u l=6.28u 
R_pattern_53 a_53 WELL ntap1 w=4.25u l=6.28u 
R_pattern_54 a_54 WELL ntap1 w=3.76u l=6.28u 
R_pattern_55 a_55 WELL ntap1 w=3.61u l=6.28u 
R_pattern_56 a_56 WELL ntap1 w=6.43u l=6.28u 
R_pattern_57 a_57 WELL ntap1 w=6.43u l=9.68u 
R_pattern_58 a_58 WELL ntap1 w=3.61u l=9.68u 
R_pattern_59 a_59 WELL ntap1 w=3.76u l=9.68u 
R_pattern_60 a_60 WELL ntap1 w=4.25u l=9.68u 
R_pattern_61 a_61 WELL ntap1 w=6.88u l=9.68u 
R_pattern_62 a_62 WELL ntap1 w=5.31u l=9.68u 
R_pattern_63 a_63 WELL ntap1 w=9.79u l=9.68u 
R_pattern_64 a_64 WELL ntap1 w=8.06u l=9.68u 
.ENDS
