VBIC Test Ic=f(Vc,Ib)

.lib ../models/cornerHBT.lib hbt_typ

ib 0 b 10u
vc c 0 1.0
vs s 0 0.0
XQ1 C B 0 S t npn13G2 nx=4

.step ib 2u 10u 2u
.dc vc 0.0 2.0 0.01
.print dc format=gnuplot v(c) i(vc) i(vs)

.end
