*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT sg13_lv_nmos
MN1 D1 G1 S1 sub sg13_lv_nmos w=150.00n l=130.00n ng=1 m=1
MN2 D2 G2 S2 digisub sg13_lv_nmos w=200.00n l=130.00n ng=1 m=1
MN3 D3 G3 S3 isosub sg13_lv_nmos w=200.00n l=150.00n ng=1 m=1
MN4 D4 G4 S4 sub sg13_lv_nmos w=300.00n l=150.00n ng=2 m=1
MN5 D5 G5 S5 sub sg13_lv_nmos w=300.00n l=300.00n ng=3 m=1
MN6 D6 G6 S6 sub sg13_lv_nmos w=200.00n l=250.00n ng=1 m=3
MN7 D7 G7 S7 sub sg13_lv_nmos w=300.00n l=150.00n ng=2 m=2

* Extra patterns
M_pattern_37 D_37 G_37 S_37 sub sg13_lv_nmos w=5.55u l=3.74u ng=1 
M_pattern_40 D_40 G_40 S_40 sub sg13_lv_nmos w=7.09u l=4.6u ng=1 
M_pattern_42 D_42 G_42 S_42 sub sg13_lv_nmos w=9.26u l=3.59u ng=1 
M_pattern_45 D_45 G_45 S_45 sub sg13_lv_nmos w=2.05u l=4.6u ng=1 
M_pattern_47 D_47 G_47 S_47 sub sg13_lv_nmos w=9.53u l=5.74u ng=1 
M_pattern_48 D_48 G_48 S_48 sub sg13_lv_nmos w=5.76u l=3.74u ng=1 
M_pattern_50 D_50 G_50 S_50 sub sg13_lv_nmos w=9.53u l=8.38u ng=1 
M_pattern_51 D_51 G_51 S_51 sub sg13_lv_nmos w=8.29u l=5.03u ng=1 
M_pattern_54 D_54 G_54 S_54 sub sg13_lv_nmos w=4.25u l=0.77u ng=1 
M_pattern_55 D_55 G_55 S_55 sub sg13_lv_nmos w=9.26u l=5.03u ng=1 
M_pattern_56 D_56 G_56 S_56 sub sg13_lv_nmos w=7.09u l=3.59u ng=1 
M_pattern_57 D_57 G_57 S_57 sub sg13_lv_nmos w=9.53u l=0.77u ng=1 
M_pattern_60 D_60 G_60 S_60 sub sg13_lv_nmos w=4.25u l=1.17u ng=1 
M_pattern_62 D_62 G_62 S_62 sub sg13_lv_nmos w=2.05u l=8.38u ng=1  
M_pattern_65 D_65 G_65 S_65 sub sg13_lv_nmos w=8.29u l=1.17u ng=1 
M_pattern_67 D_67 G_67 S_67 sub sg13_lv_nmos w=5.76u l=1.17u ng=1 
M_pattern_68 D_68 G_68 S_68 sub sg13_lv_nmos w=5.55u l=4.6u ng=1 
M_pattern_69 D_69 G_69 S_69 sub sg13_lv_nmos w=4.25u l=3.59u ng=1 
M_pattern_70 D_70 G_70 S_70 sub sg13_lv_nmos w=4.25u l=3.59u ng=1 
M_pattern_72 D_72 G_72 S_72 sub sg13_lv_nmos w=4.25u l=8.38u ng=1 
M_pattern_74 D_74 G_74 S_74 sub sg13_lv_nmos w=4.25u l=5.74u ng=1 
.ENDS
