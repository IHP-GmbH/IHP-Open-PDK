*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT pnpMPA
Q1 sub! net1 net2 pnpMPA a=1.4p   p=5.4u m=1
Q2 sub! net3 net4 pnpMPA a=1.5p   p=5.5u m=1
Q3 sub! net5 net6 pnpMPA a=1.365p p=5.3u m=1
Q4 sub! net7 net8 pnpMPA a=1.4p   p=5.4u m=3
.ENDS
