*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rfnmoshv
MN1 D1 G1 S1 B rfnmoshv w=1.0u l=0.72u ng=1 m=1
MN2 D2 G2 S2 B rfnmoshv w=2.0u l=0.72u ng=1 m=1
MN3 D3 G3 S3 B rfnmoshv w=1.0u l=1.0u  ng=1 m=1
MN4 D4 G4 S4 B rfnmoshv w=2.0u l=0.5u  ng=2 m=1
.ENDS
