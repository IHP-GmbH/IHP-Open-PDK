# ------------------------------------------------------
#
#		Copyright 2024 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Fri Jul 12 17:37:54 2024		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_4096x16_c3_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_4096x16_c3_bm_bist 0 0 ;
  SIZE 416.64 BY 618.3 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 245.01 0 245.27 0.26 ;
    END
  END A_DIN[8]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171.37 0 171.63 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 243.48 0 243.74 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 172.9 0 173.16 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.89 0 249.15 0.26 ;
    END
  END A_BM[8]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.49 0 167.75 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 250.42 0 250.68 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 165.96 0 166.22 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.755 0 250.015 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 166.625 0 166.885 0.26 ;
    END
  END A_DOUT[7]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 403.95 0 406.76 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.71 0 395.52 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 381.47 0 384.28 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.23 0 373.04 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.99 0 361.8 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.75 0 350.56 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 336.51 0 339.32 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.27 0 328.08 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.03 0 316.84 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.79 0 305.6 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 291.55 0 294.36 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.31 0 283.12 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.07 0 271.88 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 257.83 0 260.64 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.59 0 249.4 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.35 0 238.16 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.94 0 227.75 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.64 0 217.45 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 199.19 0 202 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 188.89 0 191.7 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 178.48 0 181.29 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.24 0 170.05 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156 0 158.81 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 144.76 0 147.57 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.52 0 136.33 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.28 0 125.09 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.04 0 113.85 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.8 0 102.61 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 618.3 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.57 0 412.38 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 0 401.14 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 0 389.9 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 0 378.66 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 0 367.42 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 0 356.18 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 0 344.94 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 0 333.7 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.65 0 322.46 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 308.41 0 311.22 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 297.17 0 299.98 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.93 0 288.74 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 274.69 0 277.5 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 263.45 0 266.26 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.21 0 255.02 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.97 0 243.78 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.79 0 222.6 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 209.49 0 212.3 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 204.34 0 207.15 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 194.04 0 196.85 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 0 175.67 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 0 164.43 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 0 153.19 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 0 141.95 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 0 130.71 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 0 119.47 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 0 108.23 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 0 96.99 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 30.425 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 409.57 37.065 412.38 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 37.065 401.14 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 37.065 389.9 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 37.065 378.66 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 37.065 367.42 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 37.065 356.18 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 37.065 344.94 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 37.065 333.7 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.65 37.065 322.46 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 308.41 37.065 311.22 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 297.17 37.065 299.98 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.93 37.065 288.74 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 274.69 37.065 277.5 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 263.45 37.065 266.26 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.21 37.065 255.02 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.97 37.065 243.78 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 37.065 175.67 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 37.065 164.43 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 37.065 153.19 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 37.065 141.95 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 37.065 130.71 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 37.065 119.47 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 37.065 108.23 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 37.065 96.99 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 37.065 85.75 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 37.065 74.51 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 37.065 63.27 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 37.065 52.03 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 37.065 40.79 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 37.065 29.55 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 37.065 18.31 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 37.065 7.07 618.3 ;
    END
  END VDDARRAY!
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.49 0 267.75 0.26 ;
    END
  END A_DIN[9]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 148.89 0 149.15 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 265.96 0 266.22 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.42 0 150.68 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 271.37 0 271.63 0.26 ;
    END
  END A_BM[9]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.01 0 145.27 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 272.9 0 273.16 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.48 0 143.74 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 272.235 0 272.495 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.145 0 144.405 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 289.97 0 290.23 0.26 ;
    END
  END A_DIN[10]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.41 0 126.67 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 288.44 0 288.7 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 127.94 0 128.2 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 293.85 0 294.11 0.26 ;
    END
  END A_BM[10]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.53 0 122.79 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 295.38 0 295.64 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 121 0 121.26 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.715 0 294.975 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 121.665 0 121.925 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 312.45 0 312.71 0.26 ;
    END
  END A_DIN[11]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.93 0 104.19 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 310.92 0 311.18 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 105.46 0 105.72 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 316.33 0 316.59 0.26 ;
    END
  END A_BM[11]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.05 0 100.31 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 317.86 0 318.12 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 98.52 0 98.78 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 317.195 0 317.455 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.185 0 99.445 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.93 0 335.19 0.26 ;
    END
  END A_DIN[12]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.45 0 81.71 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.4 0 333.66 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.98 0 83.24 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.81 0 339.07 0.26 ;
    END
  END A_BM[12]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.57 0 77.83 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 340.34 0 340.6 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 76.04 0 76.3 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 339.675 0 339.935 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 76.705 0 76.965 0.26 ;
    END
  END A_DOUT[3]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 357.41 0 357.67 0.26 ;
    END
  END A_DIN[13]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 58.97 0 59.23 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.88 0 356.14 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.5 0 60.76 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 361.29 0 361.55 0.26 ;
    END
  END A_BM[13]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.09 0 55.35 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 362.82 0 363.08 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 53.56 0 53.82 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 362.155 0 362.415 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.225 0 54.485 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.89 0 380.15 0.26 ;
    END
  END A_DIN[14]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.49 0 36.75 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.36 0 378.62 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 38.02 0 38.28 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 383.77 0 384.03 0.26 ;
    END
  END A_BM[14]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.61 0 32.87 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 385.3 0 385.56 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 31.08 0 31.34 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 384.635 0 384.895 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 31.745 0 32.005 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 402.37 0 402.63 0.26 ;
    END
  END A_DIN[15]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.01 0 14.27 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.84 0 401.1 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.54 0 15.8 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 406.25 0 406.51 0.26 ;
    END
  END A_BM[15]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.13 0 10.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 407.78 0 408.04 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 8.6 0 8.86 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 407.115 0 407.375 0.26 ;
    END
  END A_DOUT[15]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0345 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.265 0 9.525 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7171 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 34.349515 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.52 0 204.78 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5127 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 38.31068 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 209.11 0 209.37 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.59 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 28.783172 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 204.01 0 204.27 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3856 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 32.744337 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 208.6 0 208.86 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4519 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 33.029126 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 189.73 0 189.99 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1867 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 31.708738 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 191.26 0 191.52 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 212.17 0 212.43 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 212.68 0 212.94 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 211.15 0 211.41 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 211.66 0 211.92 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0139 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.763754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.72 0 214.98 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7487 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.443366 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.21 0 214.47 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7429 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 59.372168 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.7 0 213.96 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4777 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 58.05178 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.19 0 213.45 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.28 0 192.54 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4931 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.191934 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 192.79 0 193.05 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2323 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 51.851133 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.3 0 193.56 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9671 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.530744 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 193.81 0 194.07 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN A_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9183 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.740105 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 222.37 0 222.63 0.26 ;
    END
  END A_ADDR[9]
  PIN A_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9183 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.204381 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 222.88 0 223.14 0.26 ;
    END
  END A_BIST_ADDR[9]
  PIN A_ADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6097 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 53.730147 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.27 0 217.53 0.26 ;
    END
  END A_ADDR[10]
  PIN A_BIST_ADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 52.460543 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.78 0 218.04 0.26 ;
    END
  END A_BIST_ADDR[10]
  PIN A_ADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6359 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.902913 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.23 0 215.49 0.26 ;
    END
  END A_ADDR[11]
  PIN A_BIST_ADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6359 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.902913 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 215.74 0 216 0.26 ;
    END
  END A_BIST_ADDR[11]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8707 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.220065 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.48 0 202.74 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81105 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.923077 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.05 0 206.31 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.54 0 205.8 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8407 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.09186 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.99 0 203.25 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.874 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 12.046332 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.41 0 224.67 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8031 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 119.45135 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 17.16 LAYER Metal3 ;
      ANTENNAMAXAREACAR 1.686364 LAYER Metal2 ;
      ANTENNAMAXAREACAR 13.900125 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.03 0 205.29 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9799 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 11.079661 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 200.95 0 201.21 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9279 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.820762 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.58 0 207.84 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7211 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.812298 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 207.07 0 207.33 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7137 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.775454 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 201.46 0 201.72 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 416.64 618.3 ;
    LAYER Metal2 ;
      RECT 0.105 37.065 0.305 618.275 ;
      RECT 1.1 617.545 1.3 618.275 ;
      RECT 1.92 617.545 2.12 618.275 ;
      RECT 2.415 617.545 2.615 618.275 ;
      RECT 2.915 617.545 3.115 618.275 ;
      RECT 3.415 617.545 3.615 618.275 ;
      RECT 3.91 617.545 4.11 618.275 ;
      RECT 4.73 617.545 4.93 618.275 ;
      RECT 5.225 617.545 5.425 618.275 ;
      RECT 5.725 617.545 5.925 618.275 ;
      RECT 7.225 0.17 7.995 0.43 ;
      RECT 7.225 0.17 7.485 11.38 ;
      RECT 7.735 0.17 7.995 17.1 ;
      RECT 6.225 617.545 6.425 618.275 ;
      RECT 6.72 617.545 6.92 618.275 ;
      RECT 7.54 617.545 7.74 618.275 ;
      RECT 8.035 617.545 8.235 618.275 ;
      RECT 8.535 617.545 8.735 618.275 ;
      RECT 8.6 0.52 8.86 2.255 ;
      RECT 9.035 617.545 9.235 618.275 ;
      RECT 9.265 0.52 9.525 8.085 ;
      RECT 9.53 617.545 9.73 618.275 ;
      RECT 10.13 0.52 10.39 1.5 ;
      RECT 10.35 617.545 10.55 618.275 ;
      RECT 10.845 617.545 11.045 618.275 ;
      RECT 11.345 617.545 11.545 618.275 ;
      RECT 11.845 617.545 12.045 618.275 ;
      RECT 12.34 617.545 12.54 618.275 ;
      RECT 13.16 617.545 13.36 618.275 ;
      RECT 13.655 617.545 13.855 618.275 ;
      RECT 14.01 0.52 14.27 2.255 ;
      RECT 14.155 617.545 14.355 618.275 ;
      RECT 14.655 617.545 14.855 618.275 ;
      RECT 15.15 617.545 15.35 618.275 ;
      RECT 16.255 0.8 17.025 1.57 ;
      RECT 16.255 0.3 16.515 13.03 ;
      RECT 16.765 0.3 17.025 13.03 ;
      RECT 15.54 0.52 15.8 2.255 ;
      RECT 15.97 617.545 16.17 618.275 ;
      RECT 16.465 617.545 16.665 618.275 ;
      RECT 16.965 617.545 17.165 618.275 ;
      RECT 17.465 617.545 17.665 618.275 ;
      RECT 17.96 617.545 18.16 618.275 ;
      RECT 18.78 617.545 18.98 618.275 ;
      RECT 19.975 0.17 20.745 0.43 ;
      RECT 19.975 0.17 20.235 13.055 ;
      RECT 20.485 0.17 20.745 13.055 ;
      RECT 19.275 617.545 19.475 618.275 ;
      RECT 19.775 617.545 19.975 618.275 ;
      RECT 20.275 617.545 20.475 618.275 ;
      RECT 20.77 617.545 20.97 618.275 ;
      RECT 21.59 617.545 21.79 618.275 ;
      RECT 22.085 617.545 22.285 618.275 ;
      RECT 22.585 617.545 22.785 618.275 ;
      RECT 23.085 617.545 23.285 618.275 ;
      RECT 23.58 617.545 23.78 618.275 ;
      RECT 24.4 617.545 24.6 618.275 ;
      RECT 24.895 617.545 25.095 618.275 ;
      RECT 25.395 617.545 25.595 618.275 ;
      RECT 25.895 617.545 26.095 618.275 ;
      RECT 26.39 617.545 26.59 618.275 ;
      RECT 27.21 617.545 27.41 618.275 ;
      RECT 27.705 617.545 27.905 618.275 ;
      RECT 28.205 617.545 28.405 618.275 ;
      RECT 29.705 0.17 30.475 0.43 ;
      RECT 29.705 0.17 29.965 11.38 ;
      RECT 30.215 0.17 30.475 17.1 ;
      RECT 28.705 617.545 28.905 618.275 ;
      RECT 29.2 617.545 29.4 618.275 ;
      RECT 30.02 617.545 30.22 618.275 ;
      RECT 30.515 617.545 30.715 618.275 ;
      RECT 31.015 617.545 31.215 618.275 ;
      RECT 31.08 0.52 31.34 2.255 ;
      RECT 31.515 617.545 31.715 618.275 ;
      RECT 31.745 0.52 32.005 8.085 ;
      RECT 32.01 617.545 32.21 618.275 ;
      RECT 32.61 0.52 32.87 1.5 ;
      RECT 32.83 617.545 33.03 618.275 ;
      RECT 33.325 617.545 33.525 618.275 ;
      RECT 33.825 617.545 34.025 618.275 ;
      RECT 34.325 617.545 34.525 618.275 ;
      RECT 34.82 617.545 35.02 618.275 ;
      RECT 35.64 617.545 35.84 618.275 ;
      RECT 36.135 617.545 36.335 618.275 ;
      RECT 36.49 0.52 36.75 2.255 ;
      RECT 36.635 617.545 36.835 618.275 ;
      RECT 37.135 617.545 37.335 618.275 ;
      RECT 37.63 617.545 37.83 618.275 ;
      RECT 38.735 0.8 39.505 1.57 ;
      RECT 38.735 0.3 38.995 13.03 ;
      RECT 39.245 0.3 39.505 13.03 ;
      RECT 38.02 0.52 38.28 2.255 ;
      RECT 38.45 617.545 38.65 618.275 ;
      RECT 38.945 617.545 39.145 618.275 ;
      RECT 39.445 617.545 39.645 618.275 ;
      RECT 39.945 617.545 40.145 618.275 ;
      RECT 40.44 617.545 40.64 618.275 ;
      RECT 41.26 617.545 41.46 618.275 ;
      RECT 42.455 0.17 43.225 0.43 ;
      RECT 42.455 0.17 42.715 13.055 ;
      RECT 42.965 0.17 43.225 13.055 ;
      RECT 41.755 617.545 41.955 618.275 ;
      RECT 42.255 617.545 42.455 618.275 ;
      RECT 42.755 617.545 42.955 618.275 ;
      RECT 43.25 617.545 43.45 618.275 ;
      RECT 44.07 617.545 44.27 618.275 ;
      RECT 44.565 617.545 44.765 618.275 ;
      RECT 45.065 617.545 45.265 618.275 ;
      RECT 45.565 617.545 45.765 618.275 ;
      RECT 46.06 617.545 46.26 618.275 ;
      RECT 46.88 617.545 47.08 618.275 ;
      RECT 47.375 617.545 47.575 618.275 ;
      RECT 47.875 617.545 48.075 618.275 ;
      RECT 48.375 617.545 48.575 618.275 ;
      RECT 48.87 617.545 49.07 618.275 ;
      RECT 49.69 617.545 49.89 618.275 ;
      RECT 50.185 617.545 50.385 618.275 ;
      RECT 50.685 617.545 50.885 618.275 ;
      RECT 52.185 0.17 52.955 0.43 ;
      RECT 52.185 0.17 52.445 11.38 ;
      RECT 52.695 0.17 52.955 17.1 ;
      RECT 51.185 617.545 51.385 618.275 ;
      RECT 51.68 617.545 51.88 618.275 ;
      RECT 52.5 617.545 52.7 618.275 ;
      RECT 52.995 617.545 53.195 618.275 ;
      RECT 53.495 617.545 53.695 618.275 ;
      RECT 53.56 0.52 53.82 2.255 ;
      RECT 53.995 617.545 54.195 618.275 ;
      RECT 54.225 0.52 54.485 8.085 ;
      RECT 54.49 617.545 54.69 618.275 ;
      RECT 55.09 0.52 55.35 1.5 ;
      RECT 55.31 617.545 55.51 618.275 ;
      RECT 55.805 617.545 56.005 618.275 ;
      RECT 56.305 617.545 56.505 618.275 ;
      RECT 56.805 617.545 57.005 618.275 ;
      RECT 57.3 617.545 57.5 618.275 ;
      RECT 58.12 617.545 58.32 618.275 ;
      RECT 58.615 617.545 58.815 618.275 ;
      RECT 58.97 0.52 59.23 2.255 ;
      RECT 59.115 617.545 59.315 618.275 ;
      RECT 59.615 617.545 59.815 618.275 ;
      RECT 60.11 617.545 60.31 618.275 ;
      RECT 61.215 0.8 61.985 1.57 ;
      RECT 61.215 0.3 61.475 13.03 ;
      RECT 61.725 0.3 61.985 13.03 ;
      RECT 60.5 0.52 60.76 2.255 ;
      RECT 60.93 617.545 61.13 618.275 ;
      RECT 61.425 617.545 61.625 618.275 ;
      RECT 61.925 617.545 62.125 618.275 ;
      RECT 62.425 617.545 62.625 618.275 ;
      RECT 62.92 617.545 63.12 618.275 ;
      RECT 63.74 617.545 63.94 618.275 ;
      RECT 64.935 0.17 65.705 0.43 ;
      RECT 64.935 0.17 65.195 13.055 ;
      RECT 65.445 0.17 65.705 13.055 ;
      RECT 64.235 617.545 64.435 618.275 ;
      RECT 64.735 617.545 64.935 618.275 ;
      RECT 65.235 617.545 65.435 618.275 ;
      RECT 65.73 617.545 65.93 618.275 ;
      RECT 66.55 617.545 66.75 618.275 ;
      RECT 67.045 617.545 67.245 618.275 ;
      RECT 67.545 617.545 67.745 618.275 ;
      RECT 68.045 617.545 68.245 618.275 ;
      RECT 68.54 617.545 68.74 618.275 ;
      RECT 69.36 617.545 69.56 618.275 ;
      RECT 69.855 617.545 70.055 618.275 ;
      RECT 70.355 617.545 70.555 618.275 ;
      RECT 70.855 617.545 71.055 618.275 ;
      RECT 71.35 617.545 71.55 618.275 ;
      RECT 72.17 617.545 72.37 618.275 ;
      RECT 72.665 617.545 72.865 618.275 ;
      RECT 73.165 617.545 73.365 618.275 ;
      RECT 74.665 0.17 75.435 0.43 ;
      RECT 74.665 0.17 74.925 11.38 ;
      RECT 75.175 0.17 75.435 17.1 ;
      RECT 73.665 617.545 73.865 618.275 ;
      RECT 74.16 617.545 74.36 618.275 ;
      RECT 74.98 617.545 75.18 618.275 ;
      RECT 75.475 617.545 75.675 618.275 ;
      RECT 75.975 617.545 76.175 618.275 ;
      RECT 76.04 0.52 76.3 2.255 ;
      RECT 76.475 617.545 76.675 618.275 ;
      RECT 76.705 0.52 76.965 8.085 ;
      RECT 76.97 617.545 77.17 618.275 ;
      RECT 77.57 0.52 77.83 1.5 ;
      RECT 77.79 617.545 77.99 618.275 ;
      RECT 78.285 617.545 78.485 618.275 ;
      RECT 78.785 617.545 78.985 618.275 ;
      RECT 79.285 617.545 79.485 618.275 ;
      RECT 79.78 617.545 79.98 618.275 ;
      RECT 80.6 617.545 80.8 618.275 ;
      RECT 81.095 617.545 81.295 618.275 ;
      RECT 81.45 0.52 81.71 2.255 ;
      RECT 81.595 617.545 81.795 618.275 ;
      RECT 82.095 617.545 82.295 618.275 ;
      RECT 82.59 617.545 82.79 618.275 ;
      RECT 83.695 0.8 84.465 1.57 ;
      RECT 83.695 0.3 83.955 13.03 ;
      RECT 84.205 0.3 84.465 13.03 ;
      RECT 82.98 0.52 83.24 2.255 ;
      RECT 83.41 617.545 83.61 618.275 ;
      RECT 83.905 617.545 84.105 618.275 ;
      RECT 84.405 617.545 84.605 618.275 ;
      RECT 84.905 617.545 85.105 618.275 ;
      RECT 85.4 617.545 85.6 618.275 ;
      RECT 86.22 617.545 86.42 618.275 ;
      RECT 87.415 0.17 88.185 0.43 ;
      RECT 87.415 0.17 87.675 13.055 ;
      RECT 87.925 0.17 88.185 13.055 ;
      RECT 86.715 617.545 86.915 618.275 ;
      RECT 87.215 617.545 87.415 618.275 ;
      RECT 87.715 617.545 87.915 618.275 ;
      RECT 88.21 617.545 88.41 618.275 ;
      RECT 89.03 617.545 89.23 618.275 ;
      RECT 89.525 617.545 89.725 618.275 ;
      RECT 90.025 617.545 90.225 618.275 ;
      RECT 90.525 617.545 90.725 618.275 ;
      RECT 91.02 617.545 91.22 618.275 ;
      RECT 91.84 617.545 92.04 618.275 ;
      RECT 92.335 617.545 92.535 618.275 ;
      RECT 92.835 617.545 93.035 618.275 ;
      RECT 93.335 617.545 93.535 618.275 ;
      RECT 93.83 617.545 94.03 618.275 ;
      RECT 94.65 617.545 94.85 618.275 ;
      RECT 95.145 617.545 95.345 618.275 ;
      RECT 95.645 617.545 95.845 618.275 ;
      RECT 97.145 0.17 97.915 0.43 ;
      RECT 97.145 0.17 97.405 11.38 ;
      RECT 97.655 0.17 97.915 17.1 ;
      RECT 96.145 617.545 96.345 618.275 ;
      RECT 96.64 617.545 96.84 618.275 ;
      RECT 97.46 617.545 97.66 618.275 ;
      RECT 97.955 617.545 98.155 618.275 ;
      RECT 98.455 617.545 98.655 618.275 ;
      RECT 98.52 0.52 98.78 2.255 ;
      RECT 98.955 617.545 99.155 618.275 ;
      RECT 99.185 0.52 99.445 8.085 ;
      RECT 99.45 617.545 99.65 618.275 ;
      RECT 100.05 0.52 100.31 1.5 ;
      RECT 100.27 617.545 100.47 618.275 ;
      RECT 100.765 617.545 100.965 618.275 ;
      RECT 101.265 617.545 101.465 618.275 ;
      RECT 101.765 617.545 101.965 618.275 ;
      RECT 102.26 617.545 102.46 618.275 ;
      RECT 103.08 617.545 103.28 618.275 ;
      RECT 103.575 617.545 103.775 618.275 ;
      RECT 103.93 0.52 104.19 2.255 ;
      RECT 104.075 617.545 104.275 618.275 ;
      RECT 104.575 617.545 104.775 618.275 ;
      RECT 105.07 617.545 105.27 618.275 ;
      RECT 106.175 0.8 106.945 1.57 ;
      RECT 106.175 0.3 106.435 13.03 ;
      RECT 106.685 0.3 106.945 13.03 ;
      RECT 105.46 0.52 105.72 2.255 ;
      RECT 105.89 617.545 106.09 618.275 ;
      RECT 106.385 617.545 106.585 618.275 ;
      RECT 106.885 617.545 107.085 618.275 ;
      RECT 107.385 617.545 107.585 618.275 ;
      RECT 107.88 617.545 108.08 618.275 ;
      RECT 108.7 617.545 108.9 618.275 ;
      RECT 109.895 0.17 110.665 0.43 ;
      RECT 109.895 0.17 110.155 13.055 ;
      RECT 110.405 0.17 110.665 13.055 ;
      RECT 109.195 617.545 109.395 618.275 ;
      RECT 109.695 617.545 109.895 618.275 ;
      RECT 110.195 617.545 110.395 618.275 ;
      RECT 110.69 617.545 110.89 618.275 ;
      RECT 111.51 617.545 111.71 618.275 ;
      RECT 112.005 617.545 112.205 618.275 ;
      RECT 112.505 617.545 112.705 618.275 ;
      RECT 113.005 617.545 113.205 618.275 ;
      RECT 113.5 617.545 113.7 618.275 ;
      RECT 114.32 617.545 114.52 618.275 ;
      RECT 114.815 617.545 115.015 618.275 ;
      RECT 115.315 617.545 115.515 618.275 ;
      RECT 115.815 617.545 116.015 618.275 ;
      RECT 116.31 617.545 116.51 618.275 ;
      RECT 117.13 617.545 117.33 618.275 ;
      RECT 117.625 617.545 117.825 618.275 ;
      RECT 118.125 617.545 118.325 618.275 ;
      RECT 119.625 0.17 120.395 0.43 ;
      RECT 119.625 0.17 119.885 11.38 ;
      RECT 120.135 0.17 120.395 17.1 ;
      RECT 118.625 617.545 118.825 618.275 ;
      RECT 119.12 617.545 119.32 618.275 ;
      RECT 119.94 617.545 120.14 618.275 ;
      RECT 120.435 617.545 120.635 618.275 ;
      RECT 120.935 617.545 121.135 618.275 ;
      RECT 121 0.52 121.26 2.255 ;
      RECT 121.435 617.545 121.635 618.275 ;
      RECT 121.665 0.52 121.925 8.085 ;
      RECT 121.93 617.545 122.13 618.275 ;
      RECT 122.53 0.52 122.79 1.5 ;
      RECT 122.75 617.545 122.95 618.275 ;
      RECT 123.245 617.545 123.445 618.275 ;
      RECT 123.745 617.545 123.945 618.275 ;
      RECT 124.245 617.545 124.445 618.275 ;
      RECT 124.74 617.545 124.94 618.275 ;
      RECT 125.56 617.545 125.76 618.275 ;
      RECT 126.055 617.545 126.255 618.275 ;
      RECT 126.41 0.52 126.67 2.255 ;
      RECT 126.555 617.545 126.755 618.275 ;
      RECT 127.055 617.545 127.255 618.275 ;
      RECT 127.55 617.545 127.75 618.275 ;
      RECT 128.655 0.8 129.425 1.57 ;
      RECT 128.655 0.3 128.915 13.03 ;
      RECT 129.165 0.3 129.425 13.03 ;
      RECT 127.94 0.52 128.2 2.255 ;
      RECT 128.37 617.545 128.57 618.275 ;
      RECT 128.865 617.545 129.065 618.275 ;
      RECT 129.365 617.545 129.565 618.275 ;
      RECT 129.865 617.545 130.065 618.275 ;
      RECT 130.36 617.545 130.56 618.275 ;
      RECT 131.18 617.545 131.38 618.275 ;
      RECT 132.375 0.17 133.145 0.43 ;
      RECT 132.375 0.17 132.635 13.055 ;
      RECT 132.885 0.17 133.145 13.055 ;
      RECT 131.675 617.545 131.875 618.275 ;
      RECT 132.175 617.545 132.375 618.275 ;
      RECT 132.675 617.545 132.875 618.275 ;
      RECT 133.17 617.545 133.37 618.275 ;
      RECT 133.99 617.545 134.19 618.275 ;
      RECT 134.485 617.545 134.685 618.275 ;
      RECT 134.985 617.545 135.185 618.275 ;
      RECT 135.485 617.545 135.685 618.275 ;
      RECT 135.98 617.545 136.18 618.275 ;
      RECT 136.8 617.545 137 618.275 ;
      RECT 137.295 617.545 137.495 618.275 ;
      RECT 137.795 617.545 137.995 618.275 ;
      RECT 138.295 617.545 138.495 618.275 ;
      RECT 138.79 617.545 138.99 618.275 ;
      RECT 139.61 617.545 139.81 618.275 ;
      RECT 140.105 617.545 140.305 618.275 ;
      RECT 140.605 617.545 140.805 618.275 ;
      RECT 142.105 0.17 142.875 0.43 ;
      RECT 142.105 0.17 142.365 11.38 ;
      RECT 142.615 0.17 142.875 17.1 ;
      RECT 141.105 617.545 141.305 618.275 ;
      RECT 141.6 617.545 141.8 618.275 ;
      RECT 142.42 617.545 142.62 618.275 ;
      RECT 142.915 617.545 143.115 618.275 ;
      RECT 143.415 617.545 143.615 618.275 ;
      RECT 143.48 0.52 143.74 2.255 ;
      RECT 143.915 617.545 144.115 618.275 ;
      RECT 144.145 0.52 144.405 8.085 ;
      RECT 144.41 617.545 144.61 618.275 ;
      RECT 145.01 0.52 145.27 1.5 ;
      RECT 145.23 617.545 145.43 618.275 ;
      RECT 145.725 617.545 145.925 618.275 ;
      RECT 146.225 617.545 146.425 618.275 ;
      RECT 146.725 617.545 146.925 618.275 ;
      RECT 147.22 617.545 147.42 618.275 ;
      RECT 148.04 617.545 148.24 618.275 ;
      RECT 148.535 617.545 148.735 618.275 ;
      RECT 148.89 0.52 149.15 2.255 ;
      RECT 149.035 617.545 149.235 618.275 ;
      RECT 149.535 617.545 149.735 618.275 ;
      RECT 150.03 617.545 150.23 618.275 ;
      RECT 151.135 0.8 151.905 1.57 ;
      RECT 151.135 0.3 151.395 13.03 ;
      RECT 151.645 0.3 151.905 13.03 ;
      RECT 150.42 0.52 150.68 2.255 ;
      RECT 150.85 617.545 151.05 618.275 ;
      RECT 151.345 617.545 151.545 618.275 ;
      RECT 151.845 617.545 152.045 618.275 ;
      RECT 152.345 617.545 152.545 618.275 ;
      RECT 152.84 617.545 153.04 618.275 ;
      RECT 153.66 617.545 153.86 618.275 ;
      RECT 154.855 0.17 155.625 0.43 ;
      RECT 154.855 0.17 155.115 13.055 ;
      RECT 155.365 0.17 155.625 13.055 ;
      RECT 154.155 617.545 154.355 618.275 ;
      RECT 154.655 617.545 154.855 618.275 ;
      RECT 155.155 617.545 155.355 618.275 ;
      RECT 155.65 617.545 155.85 618.275 ;
      RECT 156.47 617.545 156.67 618.275 ;
      RECT 156.965 617.545 157.165 618.275 ;
      RECT 157.465 617.545 157.665 618.275 ;
      RECT 157.965 617.545 158.165 618.275 ;
      RECT 158.46 617.545 158.66 618.275 ;
      RECT 159.28 617.545 159.48 618.275 ;
      RECT 159.775 617.545 159.975 618.275 ;
      RECT 160.275 617.545 160.475 618.275 ;
      RECT 160.775 617.545 160.975 618.275 ;
      RECT 161.27 617.545 161.47 618.275 ;
      RECT 162.09 617.545 162.29 618.275 ;
      RECT 162.585 617.545 162.785 618.275 ;
      RECT 163.085 617.545 163.285 618.275 ;
      RECT 164.585 0.17 165.355 0.43 ;
      RECT 164.585 0.17 164.845 11.38 ;
      RECT 165.095 0.17 165.355 17.1 ;
      RECT 163.585 617.545 163.785 618.275 ;
      RECT 164.08 617.545 164.28 618.275 ;
      RECT 164.9 617.545 165.1 618.275 ;
      RECT 165.395 617.545 165.595 618.275 ;
      RECT 165.895 617.545 166.095 618.275 ;
      RECT 165.96 0.52 166.22 2.255 ;
      RECT 166.395 617.545 166.595 618.275 ;
      RECT 166.625 0.52 166.885 8.085 ;
      RECT 166.89 617.545 167.09 618.275 ;
      RECT 167.49 0.52 167.75 1.5 ;
      RECT 167.71 617.545 167.91 618.275 ;
      RECT 168.205 617.545 168.405 618.275 ;
      RECT 168.705 617.545 168.905 618.275 ;
      RECT 169.205 617.545 169.405 618.275 ;
      RECT 169.7 617.545 169.9 618.275 ;
      RECT 170.52 617.545 170.72 618.275 ;
      RECT 171.015 617.545 171.215 618.275 ;
      RECT 171.37 0.52 171.63 2.255 ;
      RECT 171.515 617.545 171.715 618.275 ;
      RECT 172.015 617.545 172.215 618.275 ;
      RECT 172.51 617.545 172.71 618.275 ;
      RECT 173.615 0.8 174.385 1.57 ;
      RECT 173.615 0.3 173.875 13.03 ;
      RECT 174.125 0.3 174.385 13.03 ;
      RECT 172.9 0.52 173.16 2.255 ;
      RECT 173.33 617.545 173.53 618.275 ;
      RECT 173.825 617.545 174.025 618.275 ;
      RECT 174.325 617.545 174.525 618.275 ;
      RECT 174.825 617.545 175.025 618.275 ;
      RECT 175.32 617.545 175.52 618.275 ;
      RECT 176.14 617.545 176.34 618.275 ;
      RECT 177.335 0.17 178.105 0.43 ;
      RECT 177.335 0.17 177.595 13.055 ;
      RECT 177.845 0.17 178.105 13.055 ;
      RECT 176.635 617.545 176.835 618.275 ;
      RECT 177.135 617.545 177.335 618.275 ;
      RECT 177.635 617.545 177.835 618.275 ;
      RECT 178.13 617.545 178.33 618.275 ;
      RECT 178.95 617.545 179.15 618.275 ;
      RECT 179.445 617.545 179.645 618.275 ;
      RECT 179.945 617.545 180.145 618.275 ;
      RECT 180.445 617.545 180.645 618.275 ;
      RECT 186.515 0.17 187.285 0.43 ;
      RECT 186.515 0.17 186.775 36.945 ;
      RECT 187.025 0.17 187.285 36.945 ;
      RECT 180.94 617.545 181.14 618.275 ;
      RECT 181.76 617.545 181.96 618.275 ;
      RECT 189.22 0 189.48 4.94 ;
      RECT 189.22 4.68 189.99 4.94 ;
      RECT 189.73 4.68 189.99 12.9 ;
      RECT 189.73 0.52 189.99 1.78 ;
      RECT 189.73 1.52 190.5 1.78 ;
      RECT 190.24 1.52 190.5 12.9 ;
      RECT 182.755 617.545 182.955 618.275 ;
      RECT 190.24 0.59 191.01 1.27 ;
      RECT 190.75 0.59 191.01 7.965 ;
      RECT 187.535 0.3 187.795 37.365 ;
      RECT 188.045 0.3 188.305 37.365 ;
      RECT 191.26 0.52 191.52 12.9 ;
      RECT 191.77 0 192.03 12.9 ;
      RECT 192.28 0.52 192.54 12.9 ;
      RECT 192.79 0.52 193.05 12.9 ;
      RECT 193.3 0.52 193.56 12.9 ;
      RECT 196.36 0.17 197.13 0.43 ;
      RECT 196.36 0.17 196.62 2.085 ;
      RECT 196.87 0.17 197.13 9 ;
      RECT 193.81 0.52 194.07 12.9 ;
      RECT 194.32 0 194.58 8.565 ;
      RECT 194.83 0 195.09 8.055 ;
      RECT 200.95 0.52 201.21 6.59 ;
      RECT 202.48 0.52 202.74 6.305 ;
      RECT 202.48 6.045 203.45 6.305 ;
      RECT 201.46 0.52 201.72 2.23 ;
      RECT 202.99 0.52 203.25 2.955 ;
      RECT 204.01 0.52 204.27 12.9 ;
      RECT 204.52 0.52 204.78 12.9 ;
      RECT 206.05 0.52 206.31 6.29 ;
      RECT 205.54 6.045 206.31 6.29 ;
      RECT 205.03 0.52 205.29 6.745 ;
      RECT 207.58 0.52 207.84 6.59 ;
      RECT 206.935 6.33 207.84 6.59 ;
      RECT 205.54 0.52 205.8 2.955 ;
      RECT 207.07 0.52 207.33 2.67 ;
      RECT 208.6 0.52 208.86 12.9 ;
      RECT 209.11 0.52 209.37 12.9 ;
      RECT 210.64 0.575 210.9 7.965 ;
      RECT 211.15 0.52 211.41 12.9 ;
      RECT 211.66 0.52 211.92 12.9 ;
      RECT 212.17 0.52 212.43 12.9 ;
      RECT 212.68 0.52 212.94 12.9 ;
      RECT 213.19 0.52 213.45 12.9 ;
      RECT 213.7 0.52 213.96 12.9 ;
      RECT 214.21 0.52 214.47 12.9 ;
      RECT 214.72 0.52 214.98 12.9 ;
      RECT 216.25 0.59 217.02 1.27 ;
      RECT 216.25 0.59 216.51 8.83 ;
      RECT 215.23 0.52 215.49 12.9 ;
      RECT 215.74 0.52 216 12.9 ;
      RECT 217.27 0.52 217.53 12.9 ;
      RECT 217.78 0.52 218.04 12.9 ;
      RECT 224.92 0.17 225.69 0.43 ;
      RECT 224.92 0.17 225.18 13.845 ;
      RECT 225.43 0.17 225.69 13.845 ;
      RECT 226.96 0.17 227.73 0.43 ;
      RECT 226.96 0.17 227.22 2.11 ;
      RECT 227.47 0.17 227.73 2.11 ;
      RECT 222.37 0.52 222.63 3.61 ;
      RECT 222.88 0.52 223.14 4.12 ;
      RECT 229.355 0.17 230.125 0.43 ;
      RECT 229.355 0.17 229.615 36.945 ;
      RECT 229.865 0.17 230.125 36.945 ;
      RECT 224.41 0.52 224.67 15.16 ;
      RECT 228.335 0.3 228.595 37.365 ;
      RECT 228.845 0.3 229.105 37.365 ;
      RECT 233.685 617.545 233.885 618.275 ;
      RECT 234.68 617.545 234.88 618.275 ;
      RECT 235.5 617.545 235.7 618.275 ;
      RECT 235.995 617.545 236.195 618.275 ;
      RECT 236.495 617.545 236.695 618.275 ;
      RECT 236.995 617.545 237.195 618.275 ;
      RECT 238.535 0.17 239.305 0.43 ;
      RECT 238.535 0.17 238.795 13.055 ;
      RECT 239.045 0.17 239.305 13.055 ;
      RECT 237.49 617.545 237.69 618.275 ;
      RECT 238.31 617.545 238.51 618.275 ;
      RECT 238.805 617.545 239.005 618.275 ;
      RECT 239.305 617.545 239.505 618.275 ;
      RECT 239.805 617.545 240.005 618.275 ;
      RECT 240.3 617.545 240.5 618.275 ;
      RECT 241.12 617.545 241.32 618.275 ;
      RECT 242.255 0.8 243.025 1.57 ;
      RECT 242.255 0.3 242.515 13.03 ;
      RECT 242.765 0.3 243.025 13.03 ;
      RECT 241.615 617.545 241.815 618.275 ;
      RECT 242.115 617.545 242.315 618.275 ;
      RECT 242.615 617.545 242.815 618.275 ;
      RECT 243.11 617.545 243.31 618.275 ;
      RECT 243.48 0.52 243.74 2.255 ;
      RECT 243.93 617.545 244.13 618.275 ;
      RECT 244.425 617.545 244.625 618.275 ;
      RECT 244.925 617.545 245.125 618.275 ;
      RECT 245.01 0.52 245.27 2.255 ;
      RECT 245.425 617.545 245.625 618.275 ;
      RECT 245.92 617.545 246.12 618.275 ;
      RECT 246.74 617.545 246.94 618.275 ;
      RECT 247.235 617.545 247.435 618.275 ;
      RECT 247.735 617.545 247.935 618.275 ;
      RECT 248.235 617.545 248.435 618.275 ;
      RECT 248.73 617.545 248.93 618.275 ;
      RECT 248.89 0.52 249.15 1.5 ;
      RECT 249.55 617.545 249.75 618.275 ;
      RECT 249.755 0.52 250.015 8.085 ;
      RECT 250.045 617.545 250.245 618.275 ;
      RECT 250.42 0.52 250.68 2.255 ;
      RECT 251.285 0.17 252.055 0.43 ;
      RECT 251.795 0.17 252.055 11.38 ;
      RECT 251.285 0.17 251.545 17.1 ;
      RECT 250.545 617.545 250.745 618.275 ;
      RECT 251.045 617.545 251.245 618.275 ;
      RECT 251.54 617.545 251.74 618.275 ;
      RECT 252.36 617.545 252.56 618.275 ;
      RECT 252.855 617.545 253.055 618.275 ;
      RECT 253.355 617.545 253.555 618.275 ;
      RECT 253.855 617.545 254.055 618.275 ;
      RECT 254.35 617.545 254.55 618.275 ;
      RECT 255.17 617.545 255.37 618.275 ;
      RECT 255.665 617.545 255.865 618.275 ;
      RECT 256.165 617.545 256.365 618.275 ;
      RECT 256.665 617.545 256.865 618.275 ;
      RECT 257.16 617.545 257.36 618.275 ;
      RECT 257.98 617.545 258.18 618.275 ;
      RECT 258.475 617.545 258.675 618.275 ;
      RECT 258.975 617.545 259.175 618.275 ;
      RECT 259.475 617.545 259.675 618.275 ;
      RECT 261.015 0.17 261.785 0.43 ;
      RECT 261.015 0.17 261.275 13.055 ;
      RECT 261.525 0.17 261.785 13.055 ;
      RECT 259.97 617.545 260.17 618.275 ;
      RECT 260.79 617.545 260.99 618.275 ;
      RECT 261.285 617.545 261.485 618.275 ;
      RECT 261.785 617.545 261.985 618.275 ;
      RECT 262.285 617.545 262.485 618.275 ;
      RECT 262.78 617.545 262.98 618.275 ;
      RECT 263.6 617.545 263.8 618.275 ;
      RECT 264.735 0.8 265.505 1.57 ;
      RECT 264.735 0.3 264.995 13.03 ;
      RECT 265.245 0.3 265.505 13.03 ;
      RECT 264.095 617.545 264.295 618.275 ;
      RECT 264.595 617.545 264.795 618.275 ;
      RECT 265.095 617.545 265.295 618.275 ;
      RECT 265.59 617.545 265.79 618.275 ;
      RECT 265.96 0.52 266.22 2.255 ;
      RECT 266.41 617.545 266.61 618.275 ;
      RECT 266.905 617.545 267.105 618.275 ;
      RECT 267.405 617.545 267.605 618.275 ;
      RECT 267.49 0.52 267.75 2.255 ;
      RECT 267.905 617.545 268.105 618.275 ;
      RECT 268.4 617.545 268.6 618.275 ;
      RECT 269.22 617.545 269.42 618.275 ;
      RECT 269.715 617.545 269.915 618.275 ;
      RECT 270.215 617.545 270.415 618.275 ;
      RECT 270.715 617.545 270.915 618.275 ;
      RECT 271.21 617.545 271.41 618.275 ;
      RECT 271.37 0.52 271.63 1.5 ;
      RECT 272.03 617.545 272.23 618.275 ;
      RECT 272.235 0.52 272.495 8.085 ;
      RECT 272.525 617.545 272.725 618.275 ;
      RECT 272.9 0.52 273.16 2.255 ;
      RECT 273.765 0.17 274.535 0.43 ;
      RECT 274.275 0.17 274.535 11.38 ;
      RECT 273.765 0.17 274.025 17.1 ;
      RECT 273.025 617.545 273.225 618.275 ;
      RECT 273.525 617.545 273.725 618.275 ;
      RECT 274.02 617.545 274.22 618.275 ;
      RECT 274.84 617.545 275.04 618.275 ;
      RECT 275.335 617.545 275.535 618.275 ;
      RECT 275.835 617.545 276.035 618.275 ;
      RECT 276.335 617.545 276.535 618.275 ;
      RECT 276.83 617.545 277.03 618.275 ;
      RECT 277.65 617.545 277.85 618.275 ;
      RECT 278.145 617.545 278.345 618.275 ;
      RECT 278.645 617.545 278.845 618.275 ;
      RECT 279.145 617.545 279.345 618.275 ;
      RECT 279.64 617.545 279.84 618.275 ;
      RECT 280.46 617.545 280.66 618.275 ;
      RECT 280.955 617.545 281.155 618.275 ;
      RECT 281.455 617.545 281.655 618.275 ;
      RECT 281.955 617.545 282.155 618.275 ;
      RECT 283.495 0.17 284.265 0.43 ;
      RECT 283.495 0.17 283.755 13.055 ;
      RECT 284.005 0.17 284.265 13.055 ;
      RECT 282.45 617.545 282.65 618.275 ;
      RECT 283.27 617.545 283.47 618.275 ;
      RECT 283.765 617.545 283.965 618.275 ;
      RECT 284.265 617.545 284.465 618.275 ;
      RECT 284.765 617.545 284.965 618.275 ;
      RECT 285.26 617.545 285.46 618.275 ;
      RECT 286.08 617.545 286.28 618.275 ;
      RECT 287.215 0.8 287.985 1.57 ;
      RECT 287.215 0.3 287.475 13.03 ;
      RECT 287.725 0.3 287.985 13.03 ;
      RECT 286.575 617.545 286.775 618.275 ;
      RECT 287.075 617.545 287.275 618.275 ;
      RECT 287.575 617.545 287.775 618.275 ;
      RECT 288.07 617.545 288.27 618.275 ;
      RECT 288.44 0.52 288.7 2.255 ;
      RECT 288.89 617.545 289.09 618.275 ;
      RECT 289.385 617.545 289.585 618.275 ;
      RECT 289.885 617.545 290.085 618.275 ;
      RECT 289.97 0.52 290.23 2.255 ;
      RECT 290.385 617.545 290.585 618.275 ;
      RECT 290.88 617.545 291.08 618.275 ;
      RECT 291.7 617.545 291.9 618.275 ;
      RECT 292.195 617.545 292.395 618.275 ;
      RECT 292.695 617.545 292.895 618.275 ;
      RECT 293.195 617.545 293.395 618.275 ;
      RECT 293.69 617.545 293.89 618.275 ;
      RECT 293.85 0.52 294.11 1.5 ;
      RECT 294.51 617.545 294.71 618.275 ;
      RECT 294.715 0.52 294.975 8.085 ;
      RECT 295.005 617.545 295.205 618.275 ;
      RECT 295.38 0.52 295.64 2.255 ;
      RECT 296.245 0.17 297.015 0.43 ;
      RECT 296.755 0.17 297.015 11.38 ;
      RECT 296.245 0.17 296.505 17.1 ;
      RECT 295.505 617.545 295.705 618.275 ;
      RECT 296.005 617.545 296.205 618.275 ;
      RECT 296.5 617.545 296.7 618.275 ;
      RECT 297.32 617.545 297.52 618.275 ;
      RECT 297.815 617.545 298.015 618.275 ;
      RECT 298.315 617.545 298.515 618.275 ;
      RECT 298.815 617.545 299.015 618.275 ;
      RECT 299.31 617.545 299.51 618.275 ;
      RECT 300.13 617.545 300.33 618.275 ;
      RECT 300.625 617.545 300.825 618.275 ;
      RECT 301.125 617.545 301.325 618.275 ;
      RECT 301.625 617.545 301.825 618.275 ;
      RECT 302.12 617.545 302.32 618.275 ;
      RECT 302.94 617.545 303.14 618.275 ;
      RECT 303.435 617.545 303.635 618.275 ;
      RECT 303.935 617.545 304.135 618.275 ;
      RECT 304.435 617.545 304.635 618.275 ;
      RECT 305.975 0.17 306.745 0.43 ;
      RECT 305.975 0.17 306.235 13.055 ;
      RECT 306.485 0.17 306.745 13.055 ;
      RECT 304.93 617.545 305.13 618.275 ;
      RECT 305.75 617.545 305.95 618.275 ;
      RECT 306.245 617.545 306.445 618.275 ;
      RECT 306.745 617.545 306.945 618.275 ;
      RECT 307.245 617.545 307.445 618.275 ;
      RECT 307.74 617.545 307.94 618.275 ;
      RECT 308.56 617.545 308.76 618.275 ;
      RECT 309.695 0.8 310.465 1.57 ;
      RECT 309.695 0.3 309.955 13.03 ;
      RECT 310.205 0.3 310.465 13.03 ;
      RECT 309.055 617.545 309.255 618.275 ;
      RECT 309.555 617.545 309.755 618.275 ;
      RECT 310.055 617.545 310.255 618.275 ;
      RECT 310.55 617.545 310.75 618.275 ;
      RECT 310.92 0.52 311.18 2.255 ;
      RECT 311.37 617.545 311.57 618.275 ;
      RECT 311.865 617.545 312.065 618.275 ;
      RECT 312.365 617.545 312.565 618.275 ;
      RECT 312.45 0.52 312.71 2.255 ;
      RECT 312.865 617.545 313.065 618.275 ;
      RECT 313.36 617.545 313.56 618.275 ;
      RECT 314.18 617.545 314.38 618.275 ;
      RECT 314.675 617.545 314.875 618.275 ;
      RECT 315.175 617.545 315.375 618.275 ;
      RECT 315.675 617.545 315.875 618.275 ;
      RECT 316.17 617.545 316.37 618.275 ;
      RECT 316.33 0.52 316.59 1.5 ;
      RECT 316.99 617.545 317.19 618.275 ;
      RECT 317.195 0.52 317.455 8.085 ;
      RECT 317.485 617.545 317.685 618.275 ;
      RECT 317.86 0.52 318.12 2.255 ;
      RECT 318.725 0.17 319.495 0.43 ;
      RECT 319.235 0.17 319.495 11.38 ;
      RECT 318.725 0.17 318.985 17.1 ;
      RECT 317.985 617.545 318.185 618.275 ;
      RECT 318.485 617.545 318.685 618.275 ;
      RECT 318.98 617.545 319.18 618.275 ;
      RECT 319.8 617.545 320 618.275 ;
      RECT 320.295 617.545 320.495 618.275 ;
      RECT 320.795 617.545 320.995 618.275 ;
      RECT 321.295 617.545 321.495 618.275 ;
      RECT 321.79 617.545 321.99 618.275 ;
      RECT 322.61 617.545 322.81 618.275 ;
      RECT 323.105 617.545 323.305 618.275 ;
      RECT 323.605 617.545 323.805 618.275 ;
      RECT 324.105 617.545 324.305 618.275 ;
      RECT 324.6 617.545 324.8 618.275 ;
      RECT 325.42 617.545 325.62 618.275 ;
      RECT 325.915 617.545 326.115 618.275 ;
      RECT 326.415 617.545 326.615 618.275 ;
      RECT 326.915 617.545 327.115 618.275 ;
      RECT 328.455 0.17 329.225 0.43 ;
      RECT 328.455 0.17 328.715 13.055 ;
      RECT 328.965 0.17 329.225 13.055 ;
      RECT 327.41 617.545 327.61 618.275 ;
      RECT 328.23 617.545 328.43 618.275 ;
      RECT 328.725 617.545 328.925 618.275 ;
      RECT 329.225 617.545 329.425 618.275 ;
      RECT 329.725 617.545 329.925 618.275 ;
      RECT 330.22 617.545 330.42 618.275 ;
      RECT 331.04 617.545 331.24 618.275 ;
      RECT 332.175 0.8 332.945 1.57 ;
      RECT 332.175 0.3 332.435 13.03 ;
      RECT 332.685 0.3 332.945 13.03 ;
      RECT 331.535 617.545 331.735 618.275 ;
      RECT 332.035 617.545 332.235 618.275 ;
      RECT 332.535 617.545 332.735 618.275 ;
      RECT 333.03 617.545 333.23 618.275 ;
      RECT 333.4 0.52 333.66 2.255 ;
      RECT 333.85 617.545 334.05 618.275 ;
      RECT 334.345 617.545 334.545 618.275 ;
      RECT 334.845 617.545 335.045 618.275 ;
      RECT 334.93 0.52 335.19 2.255 ;
      RECT 335.345 617.545 335.545 618.275 ;
      RECT 335.84 617.545 336.04 618.275 ;
      RECT 336.66 617.545 336.86 618.275 ;
      RECT 337.155 617.545 337.355 618.275 ;
      RECT 337.655 617.545 337.855 618.275 ;
      RECT 338.155 617.545 338.355 618.275 ;
      RECT 338.65 617.545 338.85 618.275 ;
      RECT 338.81 0.52 339.07 1.5 ;
      RECT 339.47 617.545 339.67 618.275 ;
      RECT 339.675 0.52 339.935 8.085 ;
      RECT 339.965 617.545 340.165 618.275 ;
      RECT 340.34 0.52 340.6 2.255 ;
      RECT 341.205 0.17 341.975 0.43 ;
      RECT 341.715 0.17 341.975 11.38 ;
      RECT 341.205 0.17 341.465 17.1 ;
      RECT 340.465 617.545 340.665 618.275 ;
      RECT 340.965 617.545 341.165 618.275 ;
      RECT 341.46 617.545 341.66 618.275 ;
      RECT 342.28 617.545 342.48 618.275 ;
      RECT 342.775 617.545 342.975 618.275 ;
      RECT 343.275 617.545 343.475 618.275 ;
      RECT 343.775 617.545 343.975 618.275 ;
      RECT 344.27 617.545 344.47 618.275 ;
      RECT 345.09 617.545 345.29 618.275 ;
      RECT 345.585 617.545 345.785 618.275 ;
      RECT 346.085 617.545 346.285 618.275 ;
      RECT 346.585 617.545 346.785 618.275 ;
      RECT 347.08 617.545 347.28 618.275 ;
      RECT 347.9 617.545 348.1 618.275 ;
      RECT 348.395 617.545 348.595 618.275 ;
      RECT 348.895 617.545 349.095 618.275 ;
      RECT 349.395 617.545 349.595 618.275 ;
      RECT 350.935 0.17 351.705 0.43 ;
      RECT 350.935 0.17 351.195 13.055 ;
      RECT 351.445 0.17 351.705 13.055 ;
      RECT 349.89 617.545 350.09 618.275 ;
      RECT 350.71 617.545 350.91 618.275 ;
      RECT 351.205 617.545 351.405 618.275 ;
      RECT 351.705 617.545 351.905 618.275 ;
      RECT 352.205 617.545 352.405 618.275 ;
      RECT 352.7 617.545 352.9 618.275 ;
      RECT 353.52 617.545 353.72 618.275 ;
      RECT 354.655 0.8 355.425 1.57 ;
      RECT 354.655 0.3 354.915 13.03 ;
      RECT 355.165 0.3 355.425 13.03 ;
      RECT 354.015 617.545 354.215 618.275 ;
      RECT 354.515 617.545 354.715 618.275 ;
      RECT 355.015 617.545 355.215 618.275 ;
      RECT 355.51 617.545 355.71 618.275 ;
      RECT 355.88 0.52 356.14 2.255 ;
      RECT 356.33 617.545 356.53 618.275 ;
      RECT 356.825 617.545 357.025 618.275 ;
      RECT 357.325 617.545 357.525 618.275 ;
      RECT 357.41 0.52 357.67 2.255 ;
      RECT 357.825 617.545 358.025 618.275 ;
      RECT 358.32 617.545 358.52 618.275 ;
      RECT 359.14 617.545 359.34 618.275 ;
      RECT 359.635 617.545 359.835 618.275 ;
      RECT 360.135 617.545 360.335 618.275 ;
      RECT 360.635 617.545 360.835 618.275 ;
      RECT 361.13 617.545 361.33 618.275 ;
      RECT 361.29 0.52 361.55 1.5 ;
      RECT 361.95 617.545 362.15 618.275 ;
      RECT 362.155 0.52 362.415 8.085 ;
      RECT 362.445 617.545 362.645 618.275 ;
      RECT 362.82 0.52 363.08 2.255 ;
      RECT 363.685 0.17 364.455 0.43 ;
      RECT 364.195 0.17 364.455 11.38 ;
      RECT 363.685 0.17 363.945 17.1 ;
      RECT 362.945 617.545 363.145 618.275 ;
      RECT 363.445 617.545 363.645 618.275 ;
      RECT 363.94 617.545 364.14 618.275 ;
      RECT 364.76 617.545 364.96 618.275 ;
      RECT 365.255 617.545 365.455 618.275 ;
      RECT 365.755 617.545 365.955 618.275 ;
      RECT 366.255 617.545 366.455 618.275 ;
      RECT 366.75 617.545 366.95 618.275 ;
      RECT 367.57 617.545 367.77 618.275 ;
      RECT 368.065 617.545 368.265 618.275 ;
      RECT 368.565 617.545 368.765 618.275 ;
      RECT 369.065 617.545 369.265 618.275 ;
      RECT 369.56 617.545 369.76 618.275 ;
      RECT 370.38 617.545 370.58 618.275 ;
      RECT 370.875 617.545 371.075 618.275 ;
      RECT 371.375 617.545 371.575 618.275 ;
      RECT 371.875 617.545 372.075 618.275 ;
      RECT 373.415 0.17 374.185 0.43 ;
      RECT 373.415 0.17 373.675 13.055 ;
      RECT 373.925 0.17 374.185 13.055 ;
      RECT 372.37 617.545 372.57 618.275 ;
      RECT 373.19 617.545 373.39 618.275 ;
      RECT 373.685 617.545 373.885 618.275 ;
      RECT 374.185 617.545 374.385 618.275 ;
      RECT 374.685 617.545 374.885 618.275 ;
      RECT 375.18 617.545 375.38 618.275 ;
      RECT 376 617.545 376.2 618.275 ;
      RECT 377.135 0.8 377.905 1.57 ;
      RECT 377.135 0.3 377.395 13.03 ;
      RECT 377.645 0.3 377.905 13.03 ;
      RECT 376.495 617.545 376.695 618.275 ;
      RECT 376.995 617.545 377.195 618.275 ;
      RECT 377.495 617.545 377.695 618.275 ;
      RECT 377.99 617.545 378.19 618.275 ;
      RECT 378.36 0.52 378.62 2.255 ;
      RECT 378.81 617.545 379.01 618.275 ;
      RECT 379.305 617.545 379.505 618.275 ;
      RECT 379.805 617.545 380.005 618.275 ;
      RECT 379.89 0.52 380.15 2.255 ;
      RECT 380.305 617.545 380.505 618.275 ;
      RECT 380.8 617.545 381 618.275 ;
      RECT 381.62 617.545 381.82 618.275 ;
      RECT 382.115 617.545 382.315 618.275 ;
      RECT 382.615 617.545 382.815 618.275 ;
      RECT 383.115 617.545 383.315 618.275 ;
      RECT 383.61 617.545 383.81 618.275 ;
      RECT 383.77 0.52 384.03 1.5 ;
      RECT 384.43 617.545 384.63 618.275 ;
      RECT 384.635 0.52 384.895 8.085 ;
      RECT 384.925 617.545 385.125 618.275 ;
      RECT 385.3 0.52 385.56 2.255 ;
      RECT 386.165 0.17 386.935 0.43 ;
      RECT 386.675 0.17 386.935 11.38 ;
      RECT 386.165 0.17 386.425 17.1 ;
      RECT 385.425 617.545 385.625 618.275 ;
      RECT 385.925 617.545 386.125 618.275 ;
      RECT 386.42 617.545 386.62 618.275 ;
      RECT 387.24 617.545 387.44 618.275 ;
      RECT 387.735 617.545 387.935 618.275 ;
      RECT 388.235 617.545 388.435 618.275 ;
      RECT 388.735 617.545 388.935 618.275 ;
      RECT 389.23 617.545 389.43 618.275 ;
      RECT 390.05 617.545 390.25 618.275 ;
      RECT 390.545 617.545 390.745 618.275 ;
      RECT 391.045 617.545 391.245 618.275 ;
      RECT 391.545 617.545 391.745 618.275 ;
      RECT 392.04 617.545 392.24 618.275 ;
      RECT 392.86 617.545 393.06 618.275 ;
      RECT 393.355 617.545 393.555 618.275 ;
      RECT 393.855 617.545 394.055 618.275 ;
      RECT 394.355 617.545 394.555 618.275 ;
      RECT 395.895 0.17 396.665 0.43 ;
      RECT 395.895 0.17 396.155 13.055 ;
      RECT 396.405 0.17 396.665 13.055 ;
      RECT 394.85 617.545 395.05 618.275 ;
      RECT 395.67 617.545 395.87 618.275 ;
      RECT 396.165 617.545 396.365 618.275 ;
      RECT 396.665 617.545 396.865 618.275 ;
      RECT 397.165 617.545 397.365 618.275 ;
      RECT 397.66 617.545 397.86 618.275 ;
      RECT 398.48 617.545 398.68 618.275 ;
      RECT 399.615 0.8 400.385 1.57 ;
      RECT 399.615 0.3 399.875 13.03 ;
      RECT 400.125 0.3 400.385 13.03 ;
      RECT 398.975 617.545 399.175 618.275 ;
      RECT 399.475 617.545 399.675 618.275 ;
      RECT 399.975 617.545 400.175 618.275 ;
      RECT 400.47 617.545 400.67 618.275 ;
      RECT 400.84 0.52 401.1 2.255 ;
      RECT 401.29 617.545 401.49 618.275 ;
      RECT 401.785 617.545 401.985 618.275 ;
      RECT 402.285 617.545 402.485 618.275 ;
      RECT 402.37 0.52 402.63 2.255 ;
      RECT 402.785 617.545 402.985 618.275 ;
      RECT 403.28 617.545 403.48 618.275 ;
      RECT 404.1 617.545 404.3 618.275 ;
      RECT 404.595 617.545 404.795 618.275 ;
      RECT 405.095 617.545 405.295 618.275 ;
      RECT 405.595 617.545 405.795 618.275 ;
      RECT 406.09 617.545 406.29 618.275 ;
      RECT 406.25 0.52 406.51 1.5 ;
      RECT 406.91 617.545 407.11 618.275 ;
      RECT 407.115 0.52 407.375 8.085 ;
      RECT 407.405 617.545 407.605 618.275 ;
      RECT 407.78 0.52 408.04 2.255 ;
      RECT 408.645 0.17 409.415 0.43 ;
      RECT 409.155 0.17 409.415 11.38 ;
      RECT 408.645 0.17 408.905 17.1 ;
      RECT 407.905 617.545 408.105 618.275 ;
      RECT 408.405 617.545 408.605 618.275 ;
      RECT 408.9 617.545 409.1 618.275 ;
      RECT 409.72 617.545 409.92 618.275 ;
      RECT 410.215 617.545 410.415 618.275 ;
      RECT 410.715 617.545 410.915 618.275 ;
      RECT 411.215 617.545 411.415 618.275 ;
      RECT 411.71 617.545 411.91 618.275 ;
      RECT 412.53 617.545 412.73 618.275 ;
      RECT 413.025 617.545 413.225 618.275 ;
      RECT 413.525 617.545 413.725 618.275 ;
      RECT 414.025 617.545 414.225 618.275 ;
      RECT 414.52 617.545 414.72 618.275 ;
      RECT 415.34 617.545 415.54 618.275 ;
      RECT 416.335 37.065 416.535 618.275 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 0 0.52 416.64 618.3 ;
      RECT 408.3 0 416.64 618.3 ;
      RECT 402.89 0 405.99 618.3 ;
      RECT 401.36 0 402.11 618.3 ;
      RECT 385.82 0 400.58 618.3 ;
      RECT 380.41 0 383.51 618.3 ;
      RECT 378.88 0 379.63 618.3 ;
      RECT 363.34 0 378.1 618.3 ;
      RECT 357.93 0 361.03 618.3 ;
      RECT 356.4 0 357.15 618.3 ;
      RECT 340.86 0 355.62 618.3 ;
      RECT 335.45 0 338.55 618.3 ;
      RECT 333.92 0 334.67 618.3 ;
      RECT 318.38 0 333.14 618.3 ;
      RECT 312.97 0 316.07 618.3 ;
      RECT 311.44 0 312.19 618.3 ;
      RECT 295.9 0 310.66 618.3 ;
      RECT 290.49 0 293.59 618.3 ;
      RECT 288.96 0 289.71 618.3 ;
      RECT 273.42 0 288.18 618.3 ;
      RECT 268.01 0 271.11 618.3 ;
      RECT 266.48 0 267.23 618.3 ;
      RECT 250.94 0 265.7 618.3 ;
      RECT 245.53 0 248.63 618.3 ;
      RECT 244 0 244.75 618.3 ;
      RECT 224.92 0.17 243.22 618.3 ;
      RECT 224.93 0 243.22 618.3 ;
      RECT 223.4 0 224.15 618.3 ;
      RECT 218.3 0 222.11 618.3 ;
      RECT 216.26 0 217.01 618.3 ;
      RECT 209.63 0 210.89 618.3 ;
      RECT 208.1 0 208.34 618.3 ;
      RECT 206.57 0 206.81 618.3 ;
      RECT 203.51 0 203.75 618.3 ;
      RECT 201.98 0 202.22 618.3 ;
      RECT 194.32 0 200.69 618.3 ;
      RECT 191.77 0 192.03 618.3 ;
      RECT 190.25 0 191 618.3 ;
      RECT 173.42 0 189.48 618.3 ;
      RECT 171.89 0 172.64 618.3 ;
      RECT 168.01 0 171.11 618.3 ;
      RECT 150.94 0 165.7 618.3 ;
      RECT 149.41 0 150.16 618.3 ;
      RECT 145.53 0 148.63 618.3 ;
      RECT 128.46 0 143.22 618.3 ;
      RECT 126.93 0 127.68 618.3 ;
      RECT 123.05 0 126.15 618.3 ;
      RECT 105.98 0 120.74 618.3 ;
      RECT 104.45 0 105.2 618.3 ;
      RECT 100.57 0 103.67 618.3 ;
      RECT 83.5 0 98.26 618.3 ;
      RECT 81.97 0 82.72 618.3 ;
      RECT 78.09 0 81.19 618.3 ;
      RECT 61.02 0 75.78 618.3 ;
      RECT 59.49 0 60.24 618.3 ;
      RECT 55.61 0 58.71 618.3 ;
      RECT 38.54 0 53.3 618.3 ;
      RECT 37.01 0 37.76 618.3 ;
      RECT 33.13 0 36.23 618.3 ;
      RECT 16.06 0 30.82 618.3 ;
      RECT 14.53 0 15.28 618.3 ;
      RECT 10.65 0 13.75 618.3 ;
      RECT 0 0 8.34 618.3 ;
    LAYER Metal3 ;
      RECT 0 0 416.64 618.3 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 228.01 0 235.09 618.3 ;
      RECT 222.86 0 224.68 618.3 ;
      RECT 217.71 0 219.53 618.3 ;
      RECT 412.64 0 416.64 618.3 ;
      RECT 407.02 0 409.31 618.3 ;
      RECT 407.02 30.685 416.64 36.805 ;
      RECT 401.4 0 403.69 618.3 ;
      RECT 395.78 0 398.07 618.3 ;
      RECT 395.78 30.685 403.69 36.805 ;
      RECT 390.16 0 392.45 618.3 ;
      RECT 384.54 0 386.83 618.3 ;
      RECT 384.54 30.685 392.45 36.805 ;
      RECT 378.92 0 381.21 618.3 ;
      RECT 373.3 0 375.59 618.3 ;
      RECT 373.3 30.685 381.21 36.805 ;
      RECT 367.68 0 369.97 618.3 ;
      RECT 362.06 0 364.35 618.3 ;
      RECT 362.06 30.685 369.97 36.805 ;
      RECT 356.44 0 358.73 618.3 ;
      RECT 350.82 0 353.11 618.3 ;
      RECT 350.82 30.685 358.73 36.805 ;
      RECT 345.2 0 347.49 618.3 ;
      RECT 339.58 0 341.87 618.3 ;
      RECT 339.58 30.685 347.49 36.805 ;
      RECT 333.96 0 336.25 618.3 ;
      RECT 328.34 0 330.63 618.3 ;
      RECT 328.34 30.685 336.25 36.805 ;
      RECT 322.72 0 325.01 618.3 ;
      RECT 317.1 0 319.39 618.3 ;
      RECT 317.1 30.685 325.01 36.805 ;
      RECT 311.48 0 313.77 618.3 ;
      RECT 305.86 0 308.15 618.3 ;
      RECT 305.86 30.685 313.77 36.805 ;
      RECT 300.24 0 302.53 618.3 ;
      RECT 80.39 0 82.68 618.3 ;
      RECT 80.39 30.685 88.3 36.805 ;
      RECT 74.77 0 77.06 618.3 ;
      RECT 69.15 0 71.44 618.3 ;
      RECT 69.15 30.685 77.06 36.805 ;
      RECT 63.53 0 65.82 618.3 ;
      RECT 57.91 0 60.2 618.3 ;
      RECT 57.91 30.685 65.82 36.805 ;
      RECT 52.29 0 54.58 618.3 ;
      RECT 46.67 0 48.96 618.3 ;
      RECT 46.67 30.685 54.58 36.805 ;
      RECT 41.05 0 43.34 618.3 ;
      RECT 35.43 0 37.72 618.3 ;
      RECT 35.43 30.685 43.34 36.805 ;
      RECT 29.81 0 32.1 618.3 ;
      RECT 24.19 0 26.48 618.3 ;
      RECT 24.19 30.685 32.1 36.805 ;
      RECT 18.57 0 20.86 618.3 ;
      RECT 12.95 0 15.24 618.3 ;
      RECT 12.95 30.685 20.86 36.805 ;
      RECT 7.33 0 9.62 618.3 ;
      RECT 0 0 4 618.3 ;
      RECT 0 30.685 9.62 36.805 ;
      RECT 294.62 0 296.91 618.3 ;
      RECT 294.62 30.685 302.53 36.805 ;
      RECT 289 0 291.29 618.3 ;
      RECT 283.38 0 285.67 618.3 ;
      RECT 283.38 30.685 291.29 36.805 ;
      RECT 277.76 0 280.05 618.3 ;
      RECT 272.14 0 274.43 618.3 ;
      RECT 272.14 30.685 280.05 36.805 ;
      RECT 266.52 0 268.81 618.3 ;
      RECT 260.9 0 263.19 618.3 ;
      RECT 260.9 30.685 268.81 36.805 ;
      RECT 255.28 0 257.57 618.3 ;
      RECT 249.66 0 251.95 618.3 ;
      RECT 249.66 30.685 257.57 36.805 ;
      RECT 244.04 0 246.33 618.3 ;
      RECT 238.42 0 240.71 618.3 ;
      RECT 238.42 30.685 246.33 36.805 ;
      RECT 212.56 0 214.38 618.3 ;
      RECT 207.41 0 209.23 618.3 ;
      RECT 202.26 0 204.08 618.3 ;
      RECT 197.11 0 198.93 618.3 ;
      RECT 191.96 0 193.78 618.3 ;
      RECT 181.55 0 188.63 618.3 ;
      RECT 175.93 0 178.22 618.3 ;
      RECT 170.31 0 172.6 618.3 ;
      RECT 170.31 30.685 178.22 36.805 ;
      RECT 164.69 0 166.98 618.3 ;
      RECT 159.07 0 161.36 618.3 ;
      RECT 159.07 30.685 166.98 36.805 ;
      RECT 153.45 0 155.74 618.3 ;
      RECT 147.83 0 150.12 618.3 ;
      RECT 147.83 30.685 155.74 36.805 ;
      RECT 142.21 0 144.5 618.3 ;
      RECT 136.59 0 138.88 618.3 ;
      RECT 136.59 30.685 144.5 36.805 ;
      RECT 130.97 0 133.26 618.3 ;
      RECT 125.35 0 127.64 618.3 ;
      RECT 125.35 30.685 133.26 36.805 ;
      RECT 119.73 0 122.02 618.3 ;
      RECT 114.11 0 116.4 618.3 ;
      RECT 114.11 30.685 122.02 36.805 ;
      RECT 108.49 0 110.78 618.3 ;
      RECT 102.87 0 105.16 618.3 ;
      RECT 102.87 30.685 110.78 36.805 ;
      RECT 97.25 0 99.54 618.3 ;
      RECT 91.63 0 93.92 618.3 ;
      RECT 91.63 30.685 99.54 36.805 ;
      RECT 86.01 0 88.3 618.3 ;
  END
END RM_IHPSG13_1P_4096x16_c3_bm_bist

END LIBRARY
