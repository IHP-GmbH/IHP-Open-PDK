########################################################################
#
# Copyright 2023 IHP PDK Authors
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#    https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
########################################################################

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_256x48_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_256x48_c2_bm_bist 0 0 ;
  SIZE 596.48 BY 118.78 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.41 0 334.67 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 261.81 0 262.07 0.26 ;
    END
  END A_DIN[23]
  PIN A_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.555 0 333.815 0.26 ;
    END
  END A_BIST_DIN[24]
  PIN A_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 262.665 0 262.925 0.26 ;
    END
  END A_BIST_DIN[23]
  PIN A_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 326.57 0 326.83 0.26 ;
    END
  END A_BM[24]
  PIN A_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 269.65 0 269.91 0.26 ;
    END
  END A_BM[23]
  PIN A_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.945 0 328.205 0.26 ;
    END
  END A_BIST_BM[24]
  PIN A_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 268.275 0 268.535 0.26 ;
    END
  END A_BIST_BM[23]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 327.08 0 327.34 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 269.14 0 269.4 0.26 ;
    END
  END A_DOUT[23]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 583.79 0 586.6 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 572.55 0 575.36 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 561.31 0 564.12 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.07 0 552.88 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 538.83 0 541.64 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 527.59 0 530.4 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 516.35 0 519.16 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 505.11 0 507.92 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 493.87 0 496.68 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 482.63 0 485.44 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 471.39 0 474.2 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 460.15 0 462.96 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.91 0 451.72 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 437.67 0 440.48 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.43 0 429.24 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 415.19 0 418 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 403.95 0 406.76 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.71 0 395.52 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 381.47 0 384.28 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.23 0 373.04 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.99 0 361.8 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.75 0 350.56 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 336.51 0 339.32 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.27 0 328.08 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 314.86 0 317.67 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 304.56 0 307.37 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 289.11 0 291.92 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278.81 0 281.62 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 268.4 0 271.21 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 257.16 0 259.97 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 245.92 0 248.73 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 234.68 0 237.49 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 223.44 0 226.25 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 212.2 0 215.01 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.96 0 203.77 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 189.72 0 192.53 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 178.48 0 181.29 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.24 0 170.05 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156 0 158.81 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 144.76 0 147.57 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.52 0 136.33 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.28 0 125.09 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.04 0 113.85 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.8 0 102.61 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.84 0 57.65 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 118.78 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 589.41 0 592.22 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.17 0 580.98 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.93 0 569.74 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.69 0 558.5 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 544.45 0 547.26 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.21 0 536.02 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 521.97 0 524.78 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 510.73 0 513.54 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 499.49 0 502.3 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.25 0 491.06 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 477.01 0 479.82 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.77 0 468.58 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 454.53 0 457.34 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 443.29 0 446.1 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 432.05 0 434.86 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 420.81 0 423.62 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.57 0 412.38 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 0 401.14 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 0 389.9 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 0 378.66 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 0 367.42 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 0 356.18 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 0 344.94 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 0 333.7 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 309.71 0 312.52 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 299.41 0 302.22 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.26 0 297.07 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 283.96 0 286.77 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.78 0 265.59 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 251.54 0 254.35 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.3 0 243.11 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 229.06 0 231.87 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.82 0 220.63 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.58 0 209.39 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.34 0 198.15 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.1 0 186.91 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 0 175.67 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 0 164.43 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 0 153.19 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 0 141.95 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 0 130.71 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 0 119.47 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 0 108.23 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 0 96.99 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 0 52.03 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 38.825 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 589.41 45.465 592.22 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 578.17 45.465 580.98 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.93 45.465 569.74 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.69 45.465 558.5 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 544.45 45.465 547.26 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.21 45.465 536.02 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 521.97 45.465 524.78 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 510.73 45.465 513.54 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 499.49 45.465 502.3 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.25 45.465 491.06 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 477.01 45.465 479.82 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.77 45.465 468.58 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 454.53 45.465 457.34 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 443.29 45.465 446.1 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 432.05 45.465 434.86 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 420.81 45.465 423.62 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.57 45.465 412.38 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 398.33 45.465 401.14 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.09 45.465 389.9 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.85 45.465 378.66 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 364.61 45.465 367.42 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 353.37 45.465 356.18 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.13 45.465 344.94 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.89 45.465 333.7 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.78 45.465 265.59 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 251.54 45.465 254.35 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.3 45.465 243.11 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 229.06 45.465 231.87 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.82 45.465 220.63 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.58 45.465 209.39 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.34 45.465 198.15 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.1 45.465 186.91 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 45.465 175.67 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 45.465 164.43 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 45.465 153.19 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 139.14 45.465 141.95 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 45.465 130.71 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 45.465 119.47 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 45.465 108.23 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.18 45.465 96.99 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 45.465 85.75 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 45.465 74.51 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 45.465 63.27 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 49.22 45.465 52.03 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 45.465 40.79 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 45.465 29.55 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 45.465 18.31 118.78 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 45.465 7.07 118.78 ;
    END
  END VDDARRAY!
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 345.65 0 345.91 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 250.57 0 250.83 0.26 ;
    END
  END A_DIN[22]
  PIN A_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 344.795 0 345.055 0.26 ;
    END
  END A_BIST_DIN[25]
  PIN A_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 251.425 0 251.685 0.26 ;
    END
  END A_BIST_DIN[22]
  PIN A_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 337.81 0 338.07 0.26 ;
    END
  END A_BM[25]
  PIN A_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 258.41 0 258.67 0.26 ;
    END
  END A_BM[22]
  PIN A_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 339.185 0 339.445 0.26 ;
    END
  END A_BIST_BM[25]
  PIN A_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 257.035 0 257.295 0.26 ;
    END
  END A_BIST_BM[22]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 338.32 0 338.58 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 257.9 0 258.16 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.89 0 357.15 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 239.33 0 239.59 0.26 ;
    END
  END A_DIN[21]
  PIN A_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.035 0 356.295 0.26 ;
    END
  END A_BIST_DIN[26]
  PIN A_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 240.185 0 240.445 0.26 ;
    END
  END A_BIST_DIN[21]
  PIN A_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.05 0 349.31 0.26 ;
    END
  END A_BM[26]
  PIN A_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 247.17 0 247.43 0.26 ;
    END
  END A_BM[21]
  PIN A_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 350.425 0 350.685 0.26 ;
    END
  END A_BIST_BM[26]
  PIN A_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 245.795 0 246.055 0.26 ;
    END
  END A_BIST_BM[21]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 349.56 0 349.82 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 246.66 0 246.92 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.13 0 368.39 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.09 0 228.35 0.26 ;
    END
  END A_DIN[20]
  PIN A_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 367.275 0 367.535 0.26 ;
    END
  END A_BIST_DIN[27]
  PIN A_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 228.945 0 229.205 0.26 ;
    END
  END A_BIST_DIN[20]
  PIN A_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.29 0 360.55 0.26 ;
    END
  END A_BM[27]
  PIN A_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 235.93 0 236.19 0.26 ;
    END
  END A_BM[20]
  PIN A_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 361.665 0 361.925 0.26 ;
    END
  END A_BIST_BM[27]
  PIN A_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 234.555 0 234.815 0.26 ;
    END
  END A_BIST_BM[20]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 360.8 0 361.06 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 235.42 0 235.68 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.37 0 379.63 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 216.85 0 217.11 0.26 ;
    END
  END A_DIN[19]
  PIN A_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 378.515 0 378.775 0.26 ;
    END
  END A_BIST_DIN[28]
  PIN A_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 217.705 0 217.965 0.26 ;
    END
  END A_BIST_DIN[19]
  PIN A_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 371.53 0 371.79 0.26 ;
    END
  END A_BM[28]
  PIN A_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.69 0 224.95 0.26 ;
    END
  END A_BM[19]
  PIN A_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.905 0 373.165 0.26 ;
    END
  END A_BIST_BM[28]
  PIN A_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 223.315 0 223.575 0.26 ;
    END
  END A_BIST_BM[19]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 372.04 0 372.3 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.18 0 224.44 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 390.61 0 390.87 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 205.61 0 205.87 0.26 ;
    END
  END A_DIN[18]
  PIN A_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 389.755 0 390.015 0.26 ;
    END
  END A_BIST_DIN[29]
  PIN A_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.465 0 206.725 0.26 ;
    END
  END A_BIST_DIN[18]
  PIN A_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 382.77 0 383.03 0.26 ;
    END
  END A_BM[29]
  PIN A_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.45 0 213.71 0.26 ;
    END
  END A_BM[18]
  PIN A_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 384.145 0 384.405 0.26 ;
    END
  END A_BIST_BM[29]
  PIN A_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 212.075 0 212.335 0.26 ;
    END
  END A_BIST_BM[18]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 383.28 0 383.54 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 212.94 0 213.2 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 401.85 0 402.11 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 194.37 0 194.63 0.26 ;
    END
  END A_DIN[17]
  PIN A_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.995 0 401.255 0.26 ;
    END
  END A_BIST_DIN[30]
  PIN A_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.225 0 195.485 0.26 ;
    END
  END A_BIST_DIN[17]
  PIN A_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 394.01 0 394.27 0.26 ;
    END
  END A_BM[30]
  PIN A_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 202.21 0 202.47 0.26 ;
    END
  END A_BM[17]
  PIN A_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 395.385 0 395.645 0.26 ;
    END
  END A_BIST_BM[30]
  PIN A_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 200.835 0 201.095 0.26 ;
    END
  END A_BIST_BM[17]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 394.52 0 394.78 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 201.7 0 201.96 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 413.09 0 413.35 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 183.13 0 183.39 0.26 ;
    END
  END A_DIN[16]
  PIN A_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 412.235 0 412.495 0.26 ;
    END
  END A_BIST_DIN[31]
  PIN A_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 183.985 0 184.245 0.26 ;
    END
  END A_BIST_DIN[16]
  PIN A_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 405.25 0 405.51 0.26 ;
    END
  END A_BM[31]
  PIN A_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 190.97 0 191.23 0.26 ;
    END
  END A_BM[16]
  PIN A_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 406.625 0 406.885 0.26 ;
    END
  END A_BIST_BM[31]
  PIN A_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 189.595 0 189.855 0.26 ;
    END
  END A_BIST_BM[16]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 405.76 0 406.02 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 190.46 0 190.72 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DIN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 424.33 0 424.59 0.26 ;
    END
  END A_DIN[32]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171.89 0 172.15 0.26 ;
    END
  END A_DIN[15]
  PIN A_BIST_DIN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 423.475 0 423.735 0.26 ;
    END
  END A_BIST_DIN[32]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 172.745 0 173.005 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BM[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 416.49 0 416.75 0.26 ;
    END
  END A_BM[32]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.73 0 179.99 0.26 ;
    END
  END A_BM[15]
  PIN A_BIST_BM[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 417.865 0 418.125 0.26 ;
    END
  END A_BIST_BM[32]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.355 0 178.615 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_DOUT[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 417 0 417.26 0.26 ;
    END
  END A_DOUT[32]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 179.22 0 179.48 0.26 ;
    END
  END A_DOUT[15]
  PIN A_DIN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 435.57 0 435.83 0.26 ;
    END
  END A_DIN[33]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.65 0 160.91 0.26 ;
    END
  END A_DIN[14]
  PIN A_BIST_DIN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 434.715 0 434.975 0.26 ;
    END
  END A_BIST_DIN[33]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.505 0 161.765 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BM[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 427.73 0 427.99 0.26 ;
    END
  END A_BM[33]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 168.49 0 168.75 0.26 ;
    END
  END A_BM[14]
  PIN A_BIST_BM[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 429.105 0 429.365 0.26 ;
    END
  END A_BIST_BM[33]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.115 0 167.375 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_DOUT[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 428.24 0 428.5 0.26 ;
    END
  END A_DOUT[33]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 167.98 0 168.24 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DIN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 446.81 0 447.07 0.26 ;
    END
  END A_DIN[34]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 149.41 0 149.67 0.26 ;
    END
  END A_DIN[13]
  PIN A_BIST_DIN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 445.955 0 446.215 0.26 ;
    END
  END A_BIST_DIN[34]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.265 0 150.525 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BM[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 438.97 0 439.23 0.26 ;
    END
  END A_BM[34]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 157.25 0 157.51 0.26 ;
    END
  END A_BM[13]
  PIN A_BIST_BM[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 440.345 0 440.605 0.26 ;
    END
  END A_BIST_BM[34]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 155.875 0 156.135 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_DOUT[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 439.48 0 439.74 0.26 ;
    END
  END A_DOUT[34]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 156.74 0 157 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DIN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 458.05 0 458.31 0.26 ;
    END
  END A_DIN[35]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 138.17 0 138.43 0.26 ;
    END
  END A_DIN[12]
  PIN A_BIST_DIN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 457.195 0 457.455 0.26 ;
    END
  END A_BIST_DIN[35]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 139.025 0 139.285 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BM[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 450.21 0 450.47 0.26 ;
    END
  END A_BM[35]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 146.01 0 146.27 0.26 ;
    END
  END A_BM[12]
  PIN A_BIST_BM[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 451.585 0 451.845 0.26 ;
    END
  END A_BIST_BM[35]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 144.635 0 144.895 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_DOUT[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 450.72 0 450.98 0.26 ;
    END
  END A_DOUT[35]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 145.5 0 145.76 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DIN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 469.29 0 469.55 0.26 ;
    END
  END A_DIN[36]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 126.93 0 127.19 0.26 ;
    END
  END A_DIN[11]
  PIN A_BIST_DIN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 468.435 0 468.695 0.26 ;
    END
  END A_BIST_DIN[36]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 127.785 0 128.045 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BM[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 461.45 0 461.71 0.26 ;
    END
  END A_BM[36]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.77 0 135.03 0.26 ;
    END
  END A_BM[11]
  PIN A_BIST_BM[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 462.825 0 463.085 0.26 ;
    END
  END A_BIST_BM[36]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.395 0 133.655 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_DOUT[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 461.96 0 462.22 0.26 ;
    END
  END A_DOUT[36]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 134.26 0 134.52 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DIN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 480.53 0 480.79 0.26 ;
    END
  END A_DIN[37]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.69 0 115.95 0.26 ;
    END
  END A_DIN[10]
  PIN A_BIST_DIN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 479.675 0 479.935 0.26 ;
    END
  END A_BIST_DIN[37]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 116.545 0 116.805 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BM[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 472.69 0 472.95 0.26 ;
    END
  END A_BM[37]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.53 0 123.79 0.26 ;
    END
  END A_BM[10]
  PIN A_BIST_BM[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 474.065 0 474.325 0.26 ;
    END
  END A_BIST_BM[37]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 122.155 0 122.415 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_DOUT[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 473.2 0 473.46 0.26 ;
    END
  END A_DOUT[37]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 123.02 0 123.28 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DIN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 491.77 0 492.03 0.26 ;
    END
  END A_DIN[38]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 104.45 0 104.71 0.26 ;
    END
  END A_DIN[9]
  PIN A_BIST_DIN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 490.915 0 491.175 0.26 ;
    END
  END A_BIST_DIN[38]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 105.305 0 105.565 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BM[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 483.93 0 484.19 0.26 ;
    END
  END A_BM[38]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 112.29 0 112.55 0.26 ;
    END
  END A_BM[9]
  PIN A_BIST_BM[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 485.305 0 485.565 0.26 ;
    END
  END A_BIST_BM[38]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 110.915 0 111.175 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_DOUT[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 484.44 0 484.7 0.26 ;
    END
  END A_DOUT[38]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 111.78 0 112.04 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DIN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 503.01 0 503.27 0.26 ;
    END
  END A_DIN[39]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 93.21 0 93.47 0.26 ;
    END
  END A_DIN[8]
  PIN A_BIST_DIN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 502.155 0 502.415 0.26 ;
    END
  END A_BIST_DIN[39]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 94.065 0 94.325 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BM[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 495.17 0 495.43 0.26 ;
    END
  END A_BM[39]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 101.05 0 101.31 0.26 ;
    END
  END A_BM[8]
  PIN A_BIST_BM[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 496.545 0 496.805 0.26 ;
    END
  END A_BIST_BM[39]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 99.675 0 99.935 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_DOUT[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 495.68 0 495.94 0.26 ;
    END
  END A_DOUT[39]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.54 0 100.8 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DIN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 514.25 0 514.51 0.26 ;
    END
  END A_DIN[40]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 81.97 0 82.23 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 513.395 0 513.655 0.26 ;
    END
  END A_BIST_DIN[40]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.825 0 83.085 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 506.41 0 506.67 0.26 ;
    END
  END A_BM[40]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.81 0 90.07 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 507.785 0 508.045 0.26 ;
    END
  END A_BIST_BM[40]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 88.435 0 88.695 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 506.92 0 507.18 0.26 ;
    END
  END A_DOUT[40]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.3 0 89.56 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DIN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 525.49 0 525.75 0.26 ;
    END
  END A_DIN[41]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.73 0 70.99 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 524.635 0 524.895 0.26 ;
    END
  END A_BIST_DIN[41]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 71.585 0 71.845 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 517.65 0 517.91 0.26 ;
    END
  END A_BM[41]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.57 0 78.83 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 519.025 0 519.285 0.26 ;
    END
  END A_BIST_BM[41]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 77.195 0 77.455 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 518.16 0 518.42 0.26 ;
    END
  END A_DOUT[41]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.06 0 78.32 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DIN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 536.73 0 536.99 0.26 ;
    END
  END A_DIN[42]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 59.49 0 59.75 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 535.875 0 536.135 0.26 ;
    END
  END A_BIST_DIN[42]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 60.345 0 60.605 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 528.89 0 529.15 0.26 ;
    END
  END A_BM[42]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 67.33 0 67.59 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 530.265 0 530.525 0.26 ;
    END
  END A_BIST_BM[42]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 65.955 0 66.215 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 529.4 0 529.66 0.26 ;
    END
  END A_DOUT[42]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 66.82 0 67.08 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DIN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 547.97 0 548.23 0.26 ;
    END
  END A_DIN[43]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 48.25 0 48.51 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 547.115 0 547.375 0.26 ;
    END
  END A_BIST_DIN[43]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 49.105 0 49.365 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 540.13 0 540.39 0.26 ;
    END
  END A_BM[43]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 56.09 0 56.35 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 541.505 0 541.765 0.26 ;
    END
  END A_BIST_BM[43]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.715 0 54.975 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 540.64 0 540.9 0.26 ;
    END
  END A_DOUT[43]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.58 0 55.84 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DIN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 559.21 0 559.47 0.26 ;
    END
  END A_DIN[44]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.01 0 37.27 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 558.355 0 558.615 0.26 ;
    END
  END A_BIST_DIN[44]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.865 0 38.125 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 551.37 0 551.63 0.26 ;
    END
  END A_BM[44]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.85 0 45.11 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 552.745 0 553.005 0.26 ;
    END
  END A_BIST_BM[44]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 43.475 0 43.735 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 551.88 0 552.14 0.26 ;
    END
  END A_DOUT[44]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.34 0 44.6 0.26 ;
    END
  END A_DOUT[3]
  PIN A_DIN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 570.45 0 570.71 0.26 ;
    END
  END A_DIN[45]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 25.77 0 26.03 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 569.595 0 569.855 0.26 ;
    END
  END A_BIST_DIN[45]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 26.625 0 26.885 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 562.61 0 562.87 0.26 ;
    END
  END A_BM[45]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.61 0 33.87 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 563.985 0 564.245 0.26 ;
    END
  END A_BIST_BM[45]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.235 0 32.495 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 563.12 0 563.38 0.26 ;
    END
  END A_DOUT[45]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.1 0 33.36 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 581.69 0 581.95 0.26 ;
    END
  END A_DIN[46]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.53 0 14.79 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 580.835 0 581.095 0.26 ;
    END
  END A_BIST_DIN[46]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.385 0 15.645 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 573.85 0 574.11 0.26 ;
    END
  END A_BM[46]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.37 0 22.63 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 575.225 0 575.485 0.26 ;
    END
  END A_BIST_BM[46]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.995 0 21.255 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 574.36 0 574.62 0.26 ;
    END
  END A_DOUT[46]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 21.86 0 22.12 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 592.93 0 593.19 0.26 ;
    END
  END A_DIN[47]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.29 0 3.55 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 592.075 0 592.335 0.26 ;
    END
  END A_BIST_DIN[47]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.145 0 4.405 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 585.09 0 585.35 0.26 ;
    END
  END A_BM[47]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.13 0 11.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 586.465 0 586.725 0.26 ;
    END
  END A_BIST_BM[47]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.755 0 10.015 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 585.6 0 585.86 0.26 ;
    END
  END A_DOUT[47]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.62 0 10.88 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 45.223301 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.44 0 294.7 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.184466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 299.03 0 299.29 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 39.656958 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 293.93 0 294.19 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.618123 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 298.52 0 298.78 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 302.09 0 302.35 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 302.6 0 302.86 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 301.07 0 301.33 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 301.58 0 301.84 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.63754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.64 0 304.9 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.317152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 304.13 0 304.39 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 70.245955 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 303.62 0 303.88 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 68.925566 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 303.11 0 303.37 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 55.436893 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 282.2 0 282.46 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 54.065721 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 282.71 0 282.97 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 62.724919 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 283.22 0 283.48 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.404531 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 283.73 0 283.99 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 292.4 0 292.66 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.796863 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 295.97 0 296.23 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 295.46 0 295.72 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 292.91 0 293.17 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 18.532819 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 314.33 0 314.59 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 292.00815 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 38.61 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.213636 LAYER Metal2 ;
      ANTENNAMAXAREACAR 17.835746 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 294.95 0 295.21 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 290.87 0 291.13 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 297.5 0 297.76 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 296.99 0 297.25 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 291.38 0 291.64 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 596.48 118.78 ;
    LAYER Metal2 ;
      RECT 0.105 45.465 0.305 118.755 ;
      RECT 1.1 118.025 1.3 118.755 ;
      RECT 3.29 0.52 3.55 5.16 ;
      RECT 2.77 4.9 3.55 5.16 ;
      RECT 2.77 4.9 3.03 6.64 ;
      RECT 1.92 118.025 2.12 118.755 ;
      RECT 2.415 118.025 2.615 118.755 ;
      RECT 2.915 118.025 3.115 118.755 ;
      RECT 3.415 118.025 3.615 118.755 ;
      RECT 3.91 118.025 4.11 118.755 ;
      RECT 4.655 0.17 5.425 0.94 ;
      RECT 4.655 0.17 4.915 12.9 ;
      RECT 5.165 0.17 5.425 12.9 ;
      RECT 4.145 0.52 4.405 5.815 ;
      RECT 4.73 118.025 4.93 118.755 ;
      RECT 5.675 0.17 6.445 0.43 ;
      RECT 5.675 0.17 5.935 11.5 ;
      RECT 6.185 0.17 6.445 11.5 ;
      RECT 5.225 118.025 5.425 118.755 ;
      RECT 5.725 118.025 5.925 118.755 ;
      RECT 6.225 118.025 6.425 118.755 ;
      RECT 7.715 0.17 8.485 0.43 ;
      RECT 7.715 0.17 7.975 10.48 ;
      RECT 8.225 0.17 8.485 10.99 ;
      RECT 6.72 118.025 6.92 118.755 ;
      RECT 7.54 118.025 7.74 118.755 ;
      RECT 8.735 0.17 9.505 0.94 ;
      RECT 8.735 0.17 8.995 8.7 ;
      RECT 9.245 0.17 9.505 12.9 ;
      RECT 8.035 118.025 8.235 118.755 ;
      RECT 8.535 118.025 8.735 118.755 ;
      RECT 9.035 118.025 9.235 118.755 ;
      RECT 9.53 118.025 9.73 118.755 ;
      RECT 9.755 0.52 10.015 2.485 ;
      RECT 10.35 118.025 10.55 118.755 ;
      RECT 10.62 0.52 10.88 14.11 ;
      RECT 10.845 118.025 11.045 118.755 ;
      RECT 11.13 0.52 11.39 2.335 ;
      RECT 11.345 118.025 11.545 118.755 ;
      RECT 11.845 118.025 12.045 118.755 ;
      RECT 12.34 118.025 12.54 118.755 ;
      RECT 14.53 0.52 14.79 5.16 ;
      RECT 14.01 4.9 14.79 5.16 ;
      RECT 14.01 4.9 14.27 6.64 ;
      RECT 13.16 118.025 13.36 118.755 ;
      RECT 13.655 118.025 13.855 118.755 ;
      RECT 14.155 118.025 14.355 118.755 ;
      RECT 14.655 118.025 14.855 118.755 ;
      RECT 15.15 118.025 15.35 118.755 ;
      RECT 15.895 0.17 16.665 0.94 ;
      RECT 15.895 0.17 16.155 12.9 ;
      RECT 16.405 0.17 16.665 12.9 ;
      RECT 15.385 0.52 15.645 5.815 ;
      RECT 15.97 118.025 16.17 118.755 ;
      RECT 16.915 0.17 17.685 0.43 ;
      RECT 16.915 0.17 17.175 11.5 ;
      RECT 17.425 0.17 17.685 11.5 ;
      RECT 16.465 118.025 16.665 118.755 ;
      RECT 16.965 118.025 17.165 118.755 ;
      RECT 17.465 118.025 17.665 118.755 ;
      RECT 18.955 0.17 19.725 0.43 ;
      RECT 18.955 0.17 19.215 10.48 ;
      RECT 19.465 0.17 19.725 10.99 ;
      RECT 17.96 118.025 18.16 118.755 ;
      RECT 18.78 118.025 18.98 118.755 ;
      RECT 19.975 0.17 20.745 0.94 ;
      RECT 19.975 0.17 20.235 8.7 ;
      RECT 20.485 0.17 20.745 12.9 ;
      RECT 19.275 118.025 19.475 118.755 ;
      RECT 19.775 118.025 19.975 118.755 ;
      RECT 20.275 118.025 20.475 118.755 ;
      RECT 20.77 118.025 20.97 118.755 ;
      RECT 20.995 0.52 21.255 2.485 ;
      RECT 21.59 118.025 21.79 118.755 ;
      RECT 21.86 0.52 22.12 14.11 ;
      RECT 22.085 118.025 22.285 118.755 ;
      RECT 22.37 0.52 22.63 2.335 ;
      RECT 22.585 118.025 22.785 118.755 ;
      RECT 23.085 118.025 23.285 118.755 ;
      RECT 23.58 118.025 23.78 118.755 ;
      RECT 25.77 0.52 26.03 5.16 ;
      RECT 25.25 4.9 26.03 5.16 ;
      RECT 25.25 4.9 25.51 6.64 ;
      RECT 24.4 118.025 24.6 118.755 ;
      RECT 24.895 118.025 25.095 118.755 ;
      RECT 25.395 118.025 25.595 118.755 ;
      RECT 25.895 118.025 26.095 118.755 ;
      RECT 26.39 118.025 26.59 118.755 ;
      RECT 27.135 0.17 27.905 0.94 ;
      RECT 27.135 0.17 27.395 12.9 ;
      RECT 27.645 0.17 27.905 12.9 ;
      RECT 26.625 0.52 26.885 5.815 ;
      RECT 27.21 118.025 27.41 118.755 ;
      RECT 28.155 0.17 28.925 0.43 ;
      RECT 28.155 0.17 28.415 11.5 ;
      RECT 28.665 0.17 28.925 11.5 ;
      RECT 27.705 118.025 27.905 118.755 ;
      RECT 28.205 118.025 28.405 118.755 ;
      RECT 28.705 118.025 28.905 118.755 ;
      RECT 30.195 0.17 30.965 0.43 ;
      RECT 30.195 0.17 30.455 10.48 ;
      RECT 30.705 0.17 30.965 10.99 ;
      RECT 29.2 118.025 29.4 118.755 ;
      RECT 30.02 118.025 30.22 118.755 ;
      RECT 31.215 0.17 31.985 0.94 ;
      RECT 31.215 0.17 31.475 8.7 ;
      RECT 31.725 0.17 31.985 12.9 ;
      RECT 30.515 118.025 30.715 118.755 ;
      RECT 31.015 118.025 31.215 118.755 ;
      RECT 31.515 118.025 31.715 118.755 ;
      RECT 32.01 118.025 32.21 118.755 ;
      RECT 32.235 0.52 32.495 2.485 ;
      RECT 32.83 118.025 33.03 118.755 ;
      RECT 33.1 0.52 33.36 14.11 ;
      RECT 33.325 118.025 33.525 118.755 ;
      RECT 33.61 0.52 33.87 2.335 ;
      RECT 33.825 118.025 34.025 118.755 ;
      RECT 34.325 118.025 34.525 118.755 ;
      RECT 34.82 118.025 35.02 118.755 ;
      RECT 37.01 0.52 37.27 5.16 ;
      RECT 36.49 4.9 37.27 5.16 ;
      RECT 36.49 4.9 36.75 6.64 ;
      RECT 35.64 118.025 35.84 118.755 ;
      RECT 36.135 118.025 36.335 118.755 ;
      RECT 36.635 118.025 36.835 118.755 ;
      RECT 37.135 118.025 37.335 118.755 ;
      RECT 37.63 118.025 37.83 118.755 ;
      RECT 38.375 0.17 39.145 0.94 ;
      RECT 38.375 0.17 38.635 12.9 ;
      RECT 38.885 0.17 39.145 12.9 ;
      RECT 37.865 0.52 38.125 5.815 ;
      RECT 38.45 118.025 38.65 118.755 ;
      RECT 39.395 0.17 40.165 0.43 ;
      RECT 39.395 0.17 39.655 11.5 ;
      RECT 39.905 0.17 40.165 11.5 ;
      RECT 38.945 118.025 39.145 118.755 ;
      RECT 39.445 118.025 39.645 118.755 ;
      RECT 39.945 118.025 40.145 118.755 ;
      RECT 41.435 0.17 42.205 0.43 ;
      RECT 41.435 0.17 41.695 10.48 ;
      RECT 41.945 0.17 42.205 10.99 ;
      RECT 40.44 118.025 40.64 118.755 ;
      RECT 41.26 118.025 41.46 118.755 ;
      RECT 42.455 0.17 43.225 0.94 ;
      RECT 42.455 0.17 42.715 8.7 ;
      RECT 42.965 0.17 43.225 12.9 ;
      RECT 41.755 118.025 41.955 118.755 ;
      RECT 42.255 118.025 42.455 118.755 ;
      RECT 42.755 118.025 42.955 118.755 ;
      RECT 43.25 118.025 43.45 118.755 ;
      RECT 43.475 0.52 43.735 2.485 ;
      RECT 44.07 118.025 44.27 118.755 ;
      RECT 44.34 0.52 44.6 14.11 ;
      RECT 44.565 118.025 44.765 118.755 ;
      RECT 44.85 0.52 45.11 2.335 ;
      RECT 45.065 118.025 45.265 118.755 ;
      RECT 45.565 118.025 45.765 118.755 ;
      RECT 46.06 118.025 46.26 118.755 ;
      RECT 48.25 0.52 48.51 5.16 ;
      RECT 47.73 4.9 48.51 5.16 ;
      RECT 47.73 4.9 47.99 6.64 ;
      RECT 46.88 118.025 47.08 118.755 ;
      RECT 47.375 118.025 47.575 118.755 ;
      RECT 47.875 118.025 48.075 118.755 ;
      RECT 48.375 118.025 48.575 118.755 ;
      RECT 48.87 118.025 49.07 118.755 ;
      RECT 49.615 0.17 50.385 0.94 ;
      RECT 49.615 0.17 49.875 12.9 ;
      RECT 50.125 0.17 50.385 12.9 ;
      RECT 49.105 0.52 49.365 5.815 ;
      RECT 49.69 118.025 49.89 118.755 ;
      RECT 50.635 0.17 51.405 0.43 ;
      RECT 50.635 0.17 50.895 11.5 ;
      RECT 51.145 0.17 51.405 11.5 ;
      RECT 50.185 118.025 50.385 118.755 ;
      RECT 50.685 118.025 50.885 118.755 ;
      RECT 51.185 118.025 51.385 118.755 ;
      RECT 52.675 0.17 53.445 0.43 ;
      RECT 52.675 0.17 52.935 10.48 ;
      RECT 53.185 0.17 53.445 10.99 ;
      RECT 51.68 118.025 51.88 118.755 ;
      RECT 52.5 118.025 52.7 118.755 ;
      RECT 53.695 0.17 54.465 0.94 ;
      RECT 53.695 0.17 53.955 8.7 ;
      RECT 54.205 0.17 54.465 12.9 ;
      RECT 52.995 118.025 53.195 118.755 ;
      RECT 53.495 118.025 53.695 118.755 ;
      RECT 53.995 118.025 54.195 118.755 ;
      RECT 54.49 118.025 54.69 118.755 ;
      RECT 54.715 0.52 54.975 2.485 ;
      RECT 55.31 118.025 55.51 118.755 ;
      RECT 55.58 0.52 55.84 14.11 ;
      RECT 55.805 118.025 56.005 118.755 ;
      RECT 56.09 0.52 56.35 2.335 ;
      RECT 56.305 118.025 56.505 118.755 ;
      RECT 56.805 118.025 57.005 118.755 ;
      RECT 57.3 118.025 57.5 118.755 ;
      RECT 59.49 0.52 59.75 5.16 ;
      RECT 58.97 4.9 59.75 5.16 ;
      RECT 58.97 4.9 59.23 6.64 ;
      RECT 58.12 118.025 58.32 118.755 ;
      RECT 58.615 118.025 58.815 118.755 ;
      RECT 59.115 118.025 59.315 118.755 ;
      RECT 59.615 118.025 59.815 118.755 ;
      RECT 60.11 118.025 60.31 118.755 ;
      RECT 60.855 0.17 61.625 0.94 ;
      RECT 60.855 0.17 61.115 12.9 ;
      RECT 61.365 0.17 61.625 12.9 ;
      RECT 60.345 0.52 60.605 5.815 ;
      RECT 60.93 118.025 61.13 118.755 ;
      RECT 61.875 0.17 62.645 0.43 ;
      RECT 61.875 0.17 62.135 11.5 ;
      RECT 62.385 0.17 62.645 11.5 ;
      RECT 61.425 118.025 61.625 118.755 ;
      RECT 61.925 118.025 62.125 118.755 ;
      RECT 62.425 118.025 62.625 118.755 ;
      RECT 63.915 0.17 64.685 0.43 ;
      RECT 63.915 0.17 64.175 10.48 ;
      RECT 64.425 0.17 64.685 10.99 ;
      RECT 62.92 118.025 63.12 118.755 ;
      RECT 63.74 118.025 63.94 118.755 ;
      RECT 64.935 0.17 65.705 0.94 ;
      RECT 64.935 0.17 65.195 8.7 ;
      RECT 65.445 0.17 65.705 12.9 ;
      RECT 64.235 118.025 64.435 118.755 ;
      RECT 64.735 118.025 64.935 118.755 ;
      RECT 65.235 118.025 65.435 118.755 ;
      RECT 65.73 118.025 65.93 118.755 ;
      RECT 65.955 0.52 66.215 2.485 ;
      RECT 66.55 118.025 66.75 118.755 ;
      RECT 66.82 0.52 67.08 14.11 ;
      RECT 67.045 118.025 67.245 118.755 ;
      RECT 67.33 0.52 67.59 2.335 ;
      RECT 67.545 118.025 67.745 118.755 ;
      RECT 68.045 118.025 68.245 118.755 ;
      RECT 68.54 118.025 68.74 118.755 ;
      RECT 70.73 0.52 70.99 5.16 ;
      RECT 70.21 4.9 70.99 5.16 ;
      RECT 70.21 4.9 70.47 6.64 ;
      RECT 69.36 118.025 69.56 118.755 ;
      RECT 69.855 118.025 70.055 118.755 ;
      RECT 70.355 118.025 70.555 118.755 ;
      RECT 70.855 118.025 71.055 118.755 ;
      RECT 71.35 118.025 71.55 118.755 ;
      RECT 72.095 0.17 72.865 0.94 ;
      RECT 72.095 0.17 72.355 12.9 ;
      RECT 72.605 0.17 72.865 12.9 ;
      RECT 71.585 0.52 71.845 5.815 ;
      RECT 72.17 118.025 72.37 118.755 ;
      RECT 73.115 0.17 73.885 0.43 ;
      RECT 73.115 0.17 73.375 11.5 ;
      RECT 73.625 0.17 73.885 11.5 ;
      RECT 72.665 118.025 72.865 118.755 ;
      RECT 73.165 118.025 73.365 118.755 ;
      RECT 73.665 118.025 73.865 118.755 ;
      RECT 75.155 0.17 75.925 0.43 ;
      RECT 75.155 0.17 75.415 10.48 ;
      RECT 75.665 0.17 75.925 10.99 ;
      RECT 74.16 118.025 74.36 118.755 ;
      RECT 74.98 118.025 75.18 118.755 ;
      RECT 76.175 0.17 76.945 0.94 ;
      RECT 76.175 0.17 76.435 8.7 ;
      RECT 76.685 0.17 76.945 12.9 ;
      RECT 75.475 118.025 75.675 118.755 ;
      RECT 75.975 118.025 76.175 118.755 ;
      RECT 76.475 118.025 76.675 118.755 ;
      RECT 76.97 118.025 77.17 118.755 ;
      RECT 77.195 0.52 77.455 2.485 ;
      RECT 77.79 118.025 77.99 118.755 ;
      RECT 78.06 0.52 78.32 14.11 ;
      RECT 78.285 118.025 78.485 118.755 ;
      RECT 78.57 0.52 78.83 2.335 ;
      RECT 78.785 118.025 78.985 118.755 ;
      RECT 79.285 118.025 79.485 118.755 ;
      RECT 79.78 118.025 79.98 118.755 ;
      RECT 81.97 0.52 82.23 5.16 ;
      RECT 81.45 4.9 82.23 5.16 ;
      RECT 81.45 4.9 81.71 6.64 ;
      RECT 80.6 118.025 80.8 118.755 ;
      RECT 81.095 118.025 81.295 118.755 ;
      RECT 81.595 118.025 81.795 118.755 ;
      RECT 82.095 118.025 82.295 118.755 ;
      RECT 82.59 118.025 82.79 118.755 ;
      RECT 83.335 0.17 84.105 0.94 ;
      RECT 83.335 0.17 83.595 12.9 ;
      RECT 83.845 0.17 84.105 12.9 ;
      RECT 82.825 0.52 83.085 5.815 ;
      RECT 83.41 118.025 83.61 118.755 ;
      RECT 84.355 0.17 85.125 0.43 ;
      RECT 84.355 0.17 84.615 11.5 ;
      RECT 84.865 0.17 85.125 11.5 ;
      RECT 83.905 118.025 84.105 118.755 ;
      RECT 84.405 118.025 84.605 118.755 ;
      RECT 84.905 118.025 85.105 118.755 ;
      RECT 86.395 0.17 87.165 0.43 ;
      RECT 86.395 0.17 86.655 10.48 ;
      RECT 86.905 0.17 87.165 10.99 ;
      RECT 85.4 118.025 85.6 118.755 ;
      RECT 86.22 118.025 86.42 118.755 ;
      RECT 87.415 0.17 88.185 0.94 ;
      RECT 87.415 0.17 87.675 8.7 ;
      RECT 87.925 0.17 88.185 12.9 ;
      RECT 86.715 118.025 86.915 118.755 ;
      RECT 87.215 118.025 87.415 118.755 ;
      RECT 87.715 118.025 87.915 118.755 ;
      RECT 88.21 118.025 88.41 118.755 ;
      RECT 88.435 0.52 88.695 2.485 ;
      RECT 89.03 118.025 89.23 118.755 ;
      RECT 89.3 0.52 89.56 14.11 ;
      RECT 89.525 118.025 89.725 118.755 ;
      RECT 89.81 0.52 90.07 2.335 ;
      RECT 90.025 118.025 90.225 118.755 ;
      RECT 90.525 118.025 90.725 118.755 ;
      RECT 91.02 118.025 91.22 118.755 ;
      RECT 93.21 0.52 93.47 5.16 ;
      RECT 92.69 4.9 93.47 5.16 ;
      RECT 92.69 4.9 92.95 6.64 ;
      RECT 91.84 118.025 92.04 118.755 ;
      RECT 92.335 118.025 92.535 118.755 ;
      RECT 92.835 118.025 93.035 118.755 ;
      RECT 93.335 118.025 93.535 118.755 ;
      RECT 93.83 118.025 94.03 118.755 ;
      RECT 94.575 0.17 95.345 0.94 ;
      RECT 94.575 0.17 94.835 12.9 ;
      RECT 95.085 0.17 95.345 12.9 ;
      RECT 94.065 0.52 94.325 5.815 ;
      RECT 94.65 118.025 94.85 118.755 ;
      RECT 95.595 0.17 96.365 0.43 ;
      RECT 95.595 0.17 95.855 11.5 ;
      RECT 96.105 0.17 96.365 11.5 ;
      RECT 95.145 118.025 95.345 118.755 ;
      RECT 95.645 118.025 95.845 118.755 ;
      RECT 96.145 118.025 96.345 118.755 ;
      RECT 97.635 0.17 98.405 0.43 ;
      RECT 97.635 0.17 97.895 10.48 ;
      RECT 98.145 0.17 98.405 10.99 ;
      RECT 96.64 118.025 96.84 118.755 ;
      RECT 97.46 118.025 97.66 118.755 ;
      RECT 98.655 0.17 99.425 0.94 ;
      RECT 98.655 0.17 98.915 8.7 ;
      RECT 99.165 0.17 99.425 12.9 ;
      RECT 97.955 118.025 98.155 118.755 ;
      RECT 98.455 118.025 98.655 118.755 ;
      RECT 98.955 118.025 99.155 118.755 ;
      RECT 99.45 118.025 99.65 118.755 ;
      RECT 99.675 0.52 99.935 2.485 ;
      RECT 100.27 118.025 100.47 118.755 ;
      RECT 100.54 0.52 100.8 14.11 ;
      RECT 100.765 118.025 100.965 118.755 ;
      RECT 101.05 0.52 101.31 2.335 ;
      RECT 101.265 118.025 101.465 118.755 ;
      RECT 101.765 118.025 101.965 118.755 ;
      RECT 102.26 118.025 102.46 118.755 ;
      RECT 104.45 0.52 104.71 5.16 ;
      RECT 103.93 4.9 104.71 5.16 ;
      RECT 103.93 4.9 104.19 6.64 ;
      RECT 103.08 118.025 103.28 118.755 ;
      RECT 103.575 118.025 103.775 118.755 ;
      RECT 104.075 118.025 104.275 118.755 ;
      RECT 104.575 118.025 104.775 118.755 ;
      RECT 105.07 118.025 105.27 118.755 ;
      RECT 105.815 0.17 106.585 0.94 ;
      RECT 105.815 0.17 106.075 12.9 ;
      RECT 106.325 0.17 106.585 12.9 ;
      RECT 105.305 0.52 105.565 5.815 ;
      RECT 105.89 118.025 106.09 118.755 ;
      RECT 106.835 0.17 107.605 0.43 ;
      RECT 106.835 0.17 107.095 11.5 ;
      RECT 107.345 0.17 107.605 11.5 ;
      RECT 106.385 118.025 106.585 118.755 ;
      RECT 106.885 118.025 107.085 118.755 ;
      RECT 107.385 118.025 107.585 118.755 ;
      RECT 108.875 0.17 109.645 0.43 ;
      RECT 108.875 0.17 109.135 10.48 ;
      RECT 109.385 0.17 109.645 10.99 ;
      RECT 107.88 118.025 108.08 118.755 ;
      RECT 108.7 118.025 108.9 118.755 ;
      RECT 109.895 0.17 110.665 0.94 ;
      RECT 109.895 0.17 110.155 8.7 ;
      RECT 110.405 0.17 110.665 12.9 ;
      RECT 109.195 118.025 109.395 118.755 ;
      RECT 109.695 118.025 109.895 118.755 ;
      RECT 110.195 118.025 110.395 118.755 ;
      RECT 110.69 118.025 110.89 118.755 ;
      RECT 110.915 0.52 111.175 2.485 ;
      RECT 111.51 118.025 111.71 118.755 ;
      RECT 111.78 0.52 112.04 14.11 ;
      RECT 112.005 118.025 112.205 118.755 ;
      RECT 112.29 0.52 112.55 2.335 ;
      RECT 112.505 118.025 112.705 118.755 ;
      RECT 113.005 118.025 113.205 118.755 ;
      RECT 113.5 118.025 113.7 118.755 ;
      RECT 115.69 0.52 115.95 5.16 ;
      RECT 115.17 4.9 115.95 5.16 ;
      RECT 115.17 4.9 115.43 6.64 ;
      RECT 114.32 118.025 114.52 118.755 ;
      RECT 114.815 118.025 115.015 118.755 ;
      RECT 115.315 118.025 115.515 118.755 ;
      RECT 115.815 118.025 116.015 118.755 ;
      RECT 116.31 118.025 116.51 118.755 ;
      RECT 117.055 0.17 117.825 0.94 ;
      RECT 117.055 0.17 117.315 12.9 ;
      RECT 117.565 0.17 117.825 12.9 ;
      RECT 116.545 0.52 116.805 5.815 ;
      RECT 117.13 118.025 117.33 118.755 ;
      RECT 118.075 0.17 118.845 0.43 ;
      RECT 118.075 0.17 118.335 11.5 ;
      RECT 118.585 0.17 118.845 11.5 ;
      RECT 117.625 118.025 117.825 118.755 ;
      RECT 118.125 118.025 118.325 118.755 ;
      RECT 118.625 118.025 118.825 118.755 ;
      RECT 120.115 0.17 120.885 0.43 ;
      RECT 120.115 0.17 120.375 10.48 ;
      RECT 120.625 0.17 120.885 10.99 ;
      RECT 119.12 118.025 119.32 118.755 ;
      RECT 119.94 118.025 120.14 118.755 ;
      RECT 121.135 0.17 121.905 0.94 ;
      RECT 121.135 0.17 121.395 8.7 ;
      RECT 121.645 0.17 121.905 12.9 ;
      RECT 120.435 118.025 120.635 118.755 ;
      RECT 120.935 118.025 121.135 118.755 ;
      RECT 121.435 118.025 121.635 118.755 ;
      RECT 121.93 118.025 122.13 118.755 ;
      RECT 122.155 0.52 122.415 2.485 ;
      RECT 122.75 118.025 122.95 118.755 ;
      RECT 123.02 0.52 123.28 14.11 ;
      RECT 123.245 118.025 123.445 118.755 ;
      RECT 123.53 0.52 123.79 2.335 ;
      RECT 123.745 118.025 123.945 118.755 ;
      RECT 124.245 118.025 124.445 118.755 ;
      RECT 124.74 118.025 124.94 118.755 ;
      RECT 126.93 0.52 127.19 5.16 ;
      RECT 126.41 4.9 127.19 5.16 ;
      RECT 126.41 4.9 126.67 6.64 ;
      RECT 125.56 118.025 125.76 118.755 ;
      RECT 126.055 118.025 126.255 118.755 ;
      RECT 126.555 118.025 126.755 118.755 ;
      RECT 127.055 118.025 127.255 118.755 ;
      RECT 127.55 118.025 127.75 118.755 ;
      RECT 128.295 0.17 129.065 0.94 ;
      RECT 128.295 0.17 128.555 12.9 ;
      RECT 128.805 0.17 129.065 12.9 ;
      RECT 127.785 0.52 128.045 5.815 ;
      RECT 128.37 118.025 128.57 118.755 ;
      RECT 129.315 0.17 130.085 0.43 ;
      RECT 129.315 0.17 129.575 11.5 ;
      RECT 129.825 0.17 130.085 11.5 ;
      RECT 128.865 118.025 129.065 118.755 ;
      RECT 129.365 118.025 129.565 118.755 ;
      RECT 129.865 118.025 130.065 118.755 ;
      RECT 131.355 0.17 132.125 0.43 ;
      RECT 131.355 0.17 131.615 10.48 ;
      RECT 131.865 0.17 132.125 10.99 ;
      RECT 130.36 118.025 130.56 118.755 ;
      RECT 131.18 118.025 131.38 118.755 ;
      RECT 132.375 0.17 133.145 0.94 ;
      RECT 132.375 0.17 132.635 8.7 ;
      RECT 132.885 0.17 133.145 12.9 ;
      RECT 131.675 118.025 131.875 118.755 ;
      RECT 132.175 118.025 132.375 118.755 ;
      RECT 132.675 118.025 132.875 118.755 ;
      RECT 133.17 118.025 133.37 118.755 ;
      RECT 133.395 0.52 133.655 2.485 ;
      RECT 133.99 118.025 134.19 118.755 ;
      RECT 134.26 0.52 134.52 14.11 ;
      RECT 134.485 118.025 134.685 118.755 ;
      RECT 134.77 0.52 135.03 2.335 ;
      RECT 134.985 118.025 135.185 118.755 ;
      RECT 135.485 118.025 135.685 118.755 ;
      RECT 135.98 118.025 136.18 118.755 ;
      RECT 138.17 0.52 138.43 5.16 ;
      RECT 137.65 4.9 138.43 5.16 ;
      RECT 137.65 4.9 137.91 6.64 ;
      RECT 136.8 118.025 137 118.755 ;
      RECT 137.295 118.025 137.495 118.755 ;
      RECT 137.795 118.025 137.995 118.755 ;
      RECT 138.295 118.025 138.495 118.755 ;
      RECT 138.79 118.025 138.99 118.755 ;
      RECT 139.535 0.17 140.305 0.94 ;
      RECT 139.535 0.17 139.795 12.9 ;
      RECT 140.045 0.17 140.305 12.9 ;
      RECT 139.025 0.52 139.285 5.815 ;
      RECT 139.61 118.025 139.81 118.755 ;
      RECT 140.555 0.17 141.325 0.43 ;
      RECT 140.555 0.17 140.815 11.5 ;
      RECT 141.065 0.17 141.325 11.5 ;
      RECT 140.105 118.025 140.305 118.755 ;
      RECT 140.605 118.025 140.805 118.755 ;
      RECT 141.105 118.025 141.305 118.755 ;
      RECT 142.595 0.17 143.365 0.43 ;
      RECT 142.595 0.17 142.855 10.48 ;
      RECT 143.105 0.17 143.365 10.99 ;
      RECT 141.6 118.025 141.8 118.755 ;
      RECT 142.42 118.025 142.62 118.755 ;
      RECT 143.615 0.17 144.385 0.94 ;
      RECT 143.615 0.17 143.875 8.7 ;
      RECT 144.125 0.17 144.385 12.9 ;
      RECT 142.915 118.025 143.115 118.755 ;
      RECT 143.415 118.025 143.615 118.755 ;
      RECT 143.915 118.025 144.115 118.755 ;
      RECT 144.41 118.025 144.61 118.755 ;
      RECT 144.635 0.52 144.895 2.485 ;
      RECT 145.23 118.025 145.43 118.755 ;
      RECT 145.5 0.52 145.76 14.11 ;
      RECT 145.725 118.025 145.925 118.755 ;
      RECT 146.01 0.52 146.27 2.335 ;
      RECT 146.225 118.025 146.425 118.755 ;
      RECT 146.725 118.025 146.925 118.755 ;
      RECT 147.22 118.025 147.42 118.755 ;
      RECT 149.41 0.52 149.67 5.16 ;
      RECT 148.89 4.9 149.67 5.16 ;
      RECT 148.89 4.9 149.15 6.64 ;
      RECT 148.04 118.025 148.24 118.755 ;
      RECT 148.535 118.025 148.735 118.755 ;
      RECT 149.035 118.025 149.235 118.755 ;
      RECT 149.535 118.025 149.735 118.755 ;
      RECT 150.03 118.025 150.23 118.755 ;
      RECT 150.775 0.17 151.545 0.94 ;
      RECT 150.775 0.17 151.035 12.9 ;
      RECT 151.285 0.17 151.545 12.9 ;
      RECT 150.265 0.52 150.525 5.815 ;
      RECT 150.85 118.025 151.05 118.755 ;
      RECT 151.795 0.17 152.565 0.43 ;
      RECT 151.795 0.17 152.055 11.5 ;
      RECT 152.305 0.17 152.565 11.5 ;
      RECT 151.345 118.025 151.545 118.755 ;
      RECT 151.845 118.025 152.045 118.755 ;
      RECT 152.345 118.025 152.545 118.755 ;
      RECT 153.835 0.17 154.605 0.43 ;
      RECT 153.835 0.17 154.095 10.48 ;
      RECT 154.345 0.17 154.605 10.99 ;
      RECT 152.84 118.025 153.04 118.755 ;
      RECT 153.66 118.025 153.86 118.755 ;
      RECT 154.855 0.17 155.625 0.94 ;
      RECT 154.855 0.17 155.115 8.7 ;
      RECT 155.365 0.17 155.625 12.9 ;
      RECT 154.155 118.025 154.355 118.755 ;
      RECT 154.655 118.025 154.855 118.755 ;
      RECT 155.155 118.025 155.355 118.755 ;
      RECT 155.65 118.025 155.85 118.755 ;
      RECT 155.875 0.52 156.135 2.485 ;
      RECT 156.47 118.025 156.67 118.755 ;
      RECT 156.74 0.52 157 14.11 ;
      RECT 156.965 118.025 157.165 118.755 ;
      RECT 157.25 0.52 157.51 2.335 ;
      RECT 157.465 118.025 157.665 118.755 ;
      RECT 157.965 118.025 158.165 118.755 ;
      RECT 158.46 118.025 158.66 118.755 ;
      RECT 160.65 0.52 160.91 5.16 ;
      RECT 160.13 4.9 160.91 5.16 ;
      RECT 160.13 4.9 160.39 6.64 ;
      RECT 159.28 118.025 159.48 118.755 ;
      RECT 159.775 118.025 159.975 118.755 ;
      RECT 160.275 118.025 160.475 118.755 ;
      RECT 160.775 118.025 160.975 118.755 ;
      RECT 161.27 118.025 161.47 118.755 ;
      RECT 162.015 0.17 162.785 0.94 ;
      RECT 162.015 0.17 162.275 12.9 ;
      RECT 162.525 0.17 162.785 12.9 ;
      RECT 161.505 0.52 161.765 5.815 ;
      RECT 162.09 118.025 162.29 118.755 ;
      RECT 163.035 0.17 163.805 0.43 ;
      RECT 163.035 0.17 163.295 11.5 ;
      RECT 163.545 0.17 163.805 11.5 ;
      RECT 162.585 118.025 162.785 118.755 ;
      RECT 163.085 118.025 163.285 118.755 ;
      RECT 163.585 118.025 163.785 118.755 ;
      RECT 165.075 0.17 165.845 0.43 ;
      RECT 165.075 0.17 165.335 10.48 ;
      RECT 165.585 0.17 165.845 10.99 ;
      RECT 164.08 118.025 164.28 118.755 ;
      RECT 164.9 118.025 165.1 118.755 ;
      RECT 166.095 0.17 166.865 0.94 ;
      RECT 166.095 0.17 166.355 8.7 ;
      RECT 166.605 0.17 166.865 12.9 ;
      RECT 165.395 118.025 165.595 118.755 ;
      RECT 165.895 118.025 166.095 118.755 ;
      RECT 166.395 118.025 166.595 118.755 ;
      RECT 166.89 118.025 167.09 118.755 ;
      RECT 167.115 0.52 167.375 2.485 ;
      RECT 167.71 118.025 167.91 118.755 ;
      RECT 167.98 0.52 168.24 14.11 ;
      RECT 168.205 118.025 168.405 118.755 ;
      RECT 168.49 0.52 168.75 2.335 ;
      RECT 168.705 118.025 168.905 118.755 ;
      RECT 169.205 118.025 169.405 118.755 ;
      RECT 169.7 118.025 169.9 118.755 ;
      RECT 171.89 0.52 172.15 5.16 ;
      RECT 171.37 4.9 172.15 5.16 ;
      RECT 171.37 4.9 171.63 6.64 ;
      RECT 170.52 118.025 170.72 118.755 ;
      RECT 171.015 118.025 171.215 118.755 ;
      RECT 171.515 118.025 171.715 118.755 ;
      RECT 172.015 118.025 172.215 118.755 ;
      RECT 172.51 118.025 172.71 118.755 ;
      RECT 173.255 0.17 174.025 0.94 ;
      RECT 173.255 0.17 173.515 12.9 ;
      RECT 173.765 0.17 174.025 12.9 ;
      RECT 172.745 0.52 173.005 5.815 ;
      RECT 173.33 118.025 173.53 118.755 ;
      RECT 174.275 0.17 175.045 0.43 ;
      RECT 174.275 0.17 174.535 11.5 ;
      RECT 174.785 0.17 175.045 11.5 ;
      RECT 173.825 118.025 174.025 118.755 ;
      RECT 174.325 118.025 174.525 118.755 ;
      RECT 174.825 118.025 175.025 118.755 ;
      RECT 176.315 0.17 177.085 0.43 ;
      RECT 176.315 0.17 176.575 10.48 ;
      RECT 176.825 0.17 177.085 10.99 ;
      RECT 175.32 118.025 175.52 118.755 ;
      RECT 176.14 118.025 176.34 118.755 ;
      RECT 177.335 0.17 178.105 0.94 ;
      RECT 177.335 0.17 177.595 8.7 ;
      RECT 177.845 0.17 178.105 12.9 ;
      RECT 176.635 118.025 176.835 118.755 ;
      RECT 177.135 118.025 177.335 118.755 ;
      RECT 177.635 118.025 177.835 118.755 ;
      RECT 178.13 118.025 178.33 118.755 ;
      RECT 178.355 0.52 178.615 2.485 ;
      RECT 178.95 118.025 179.15 118.755 ;
      RECT 179.22 0.52 179.48 14.11 ;
      RECT 179.445 118.025 179.645 118.755 ;
      RECT 179.73 0.52 179.99 2.335 ;
      RECT 179.945 118.025 180.145 118.755 ;
      RECT 180.445 118.025 180.645 118.755 ;
      RECT 180.94 118.025 181.14 118.755 ;
      RECT 183.13 0.52 183.39 5.16 ;
      RECT 182.61 4.9 183.39 5.16 ;
      RECT 182.61 4.9 182.87 6.64 ;
      RECT 181.76 118.025 181.96 118.755 ;
      RECT 182.255 118.025 182.455 118.755 ;
      RECT 182.755 118.025 182.955 118.755 ;
      RECT 183.255 118.025 183.455 118.755 ;
      RECT 183.75 118.025 183.95 118.755 ;
      RECT 184.495 0.17 185.265 0.94 ;
      RECT 184.495 0.17 184.755 12.9 ;
      RECT 185.005 0.17 185.265 12.9 ;
      RECT 183.985 0.52 184.245 5.815 ;
      RECT 184.57 118.025 184.77 118.755 ;
      RECT 185.515 0.17 186.285 0.43 ;
      RECT 185.515 0.17 185.775 11.5 ;
      RECT 186.025 0.17 186.285 11.5 ;
      RECT 185.065 118.025 185.265 118.755 ;
      RECT 185.565 118.025 185.765 118.755 ;
      RECT 186.065 118.025 186.265 118.755 ;
      RECT 187.555 0.17 188.325 0.43 ;
      RECT 187.555 0.17 187.815 10.48 ;
      RECT 188.065 0.17 188.325 10.99 ;
      RECT 186.56 118.025 186.76 118.755 ;
      RECT 187.38 118.025 187.58 118.755 ;
      RECT 188.575 0.17 189.345 0.94 ;
      RECT 188.575 0.17 188.835 8.7 ;
      RECT 189.085 0.17 189.345 12.9 ;
      RECT 187.875 118.025 188.075 118.755 ;
      RECT 188.375 118.025 188.575 118.755 ;
      RECT 188.875 118.025 189.075 118.755 ;
      RECT 189.37 118.025 189.57 118.755 ;
      RECT 189.595 0.52 189.855 2.485 ;
      RECT 190.19 118.025 190.39 118.755 ;
      RECT 190.46 0.52 190.72 14.11 ;
      RECT 190.685 118.025 190.885 118.755 ;
      RECT 190.97 0.52 191.23 2.335 ;
      RECT 191.185 118.025 191.385 118.755 ;
      RECT 191.685 118.025 191.885 118.755 ;
      RECT 192.18 118.025 192.38 118.755 ;
      RECT 194.37 0.52 194.63 5.16 ;
      RECT 193.85 4.9 194.63 5.16 ;
      RECT 193.85 4.9 194.11 6.64 ;
      RECT 193 118.025 193.2 118.755 ;
      RECT 193.495 118.025 193.695 118.755 ;
      RECT 193.995 118.025 194.195 118.755 ;
      RECT 194.495 118.025 194.695 118.755 ;
      RECT 194.99 118.025 195.19 118.755 ;
      RECT 195.735 0.17 196.505 0.94 ;
      RECT 195.735 0.17 195.995 12.9 ;
      RECT 196.245 0.17 196.505 12.9 ;
      RECT 195.225 0.52 195.485 5.815 ;
      RECT 195.81 118.025 196.01 118.755 ;
      RECT 196.755 0.17 197.525 0.43 ;
      RECT 196.755 0.17 197.015 11.5 ;
      RECT 197.265 0.17 197.525 11.5 ;
      RECT 196.305 118.025 196.505 118.755 ;
      RECT 196.805 118.025 197.005 118.755 ;
      RECT 197.305 118.025 197.505 118.755 ;
      RECT 198.795 0.17 199.565 0.43 ;
      RECT 198.795 0.17 199.055 10.48 ;
      RECT 199.305 0.17 199.565 10.99 ;
      RECT 197.8 118.025 198 118.755 ;
      RECT 198.62 118.025 198.82 118.755 ;
      RECT 199.815 0.17 200.585 0.94 ;
      RECT 199.815 0.17 200.075 8.7 ;
      RECT 200.325 0.17 200.585 12.9 ;
      RECT 199.115 118.025 199.315 118.755 ;
      RECT 199.615 118.025 199.815 118.755 ;
      RECT 200.115 118.025 200.315 118.755 ;
      RECT 200.61 118.025 200.81 118.755 ;
      RECT 200.835 0.52 201.095 2.485 ;
      RECT 201.43 118.025 201.63 118.755 ;
      RECT 201.7 0.52 201.96 14.11 ;
      RECT 201.925 118.025 202.125 118.755 ;
      RECT 202.21 0.52 202.47 2.335 ;
      RECT 202.425 118.025 202.625 118.755 ;
      RECT 202.925 118.025 203.125 118.755 ;
      RECT 203.42 118.025 203.62 118.755 ;
      RECT 205.61 0.52 205.87 5.16 ;
      RECT 205.09 4.9 205.87 5.16 ;
      RECT 205.09 4.9 205.35 6.64 ;
      RECT 204.24 118.025 204.44 118.755 ;
      RECT 204.735 118.025 204.935 118.755 ;
      RECT 205.235 118.025 205.435 118.755 ;
      RECT 205.735 118.025 205.935 118.755 ;
      RECT 206.23 118.025 206.43 118.755 ;
      RECT 206.975 0.17 207.745 0.94 ;
      RECT 206.975 0.17 207.235 12.9 ;
      RECT 207.485 0.17 207.745 12.9 ;
      RECT 206.465 0.52 206.725 5.815 ;
      RECT 207.05 118.025 207.25 118.755 ;
      RECT 207.995 0.17 208.765 0.43 ;
      RECT 207.995 0.17 208.255 11.5 ;
      RECT 208.505 0.17 208.765 11.5 ;
      RECT 207.545 118.025 207.745 118.755 ;
      RECT 208.045 118.025 208.245 118.755 ;
      RECT 208.545 118.025 208.745 118.755 ;
      RECT 210.035 0.17 210.805 0.43 ;
      RECT 210.035 0.17 210.295 10.48 ;
      RECT 210.545 0.17 210.805 10.99 ;
      RECT 209.04 118.025 209.24 118.755 ;
      RECT 209.86 118.025 210.06 118.755 ;
      RECT 211.055 0.17 211.825 0.94 ;
      RECT 211.055 0.17 211.315 8.7 ;
      RECT 211.565 0.17 211.825 12.9 ;
      RECT 210.355 118.025 210.555 118.755 ;
      RECT 210.855 118.025 211.055 118.755 ;
      RECT 211.355 118.025 211.555 118.755 ;
      RECT 211.85 118.025 212.05 118.755 ;
      RECT 212.075 0.52 212.335 2.485 ;
      RECT 212.67 118.025 212.87 118.755 ;
      RECT 212.94 0.52 213.2 14.11 ;
      RECT 213.165 118.025 213.365 118.755 ;
      RECT 213.45 0.52 213.71 2.335 ;
      RECT 213.665 118.025 213.865 118.755 ;
      RECT 214.165 118.025 214.365 118.755 ;
      RECT 214.66 118.025 214.86 118.755 ;
      RECT 216.85 0.52 217.11 5.16 ;
      RECT 216.33 4.9 217.11 5.16 ;
      RECT 216.33 4.9 216.59 6.64 ;
      RECT 215.48 118.025 215.68 118.755 ;
      RECT 215.975 118.025 216.175 118.755 ;
      RECT 216.475 118.025 216.675 118.755 ;
      RECT 216.975 118.025 217.175 118.755 ;
      RECT 217.47 118.025 217.67 118.755 ;
      RECT 218.215 0.17 218.985 0.94 ;
      RECT 218.215 0.17 218.475 12.9 ;
      RECT 218.725 0.17 218.985 12.9 ;
      RECT 217.705 0.52 217.965 5.815 ;
      RECT 218.29 118.025 218.49 118.755 ;
      RECT 219.235 0.17 220.005 0.43 ;
      RECT 219.235 0.17 219.495 11.5 ;
      RECT 219.745 0.17 220.005 11.5 ;
      RECT 218.785 118.025 218.985 118.755 ;
      RECT 219.285 118.025 219.485 118.755 ;
      RECT 219.785 118.025 219.985 118.755 ;
      RECT 221.275 0.17 222.045 0.43 ;
      RECT 221.275 0.17 221.535 10.48 ;
      RECT 221.785 0.17 222.045 10.99 ;
      RECT 220.28 118.025 220.48 118.755 ;
      RECT 221.1 118.025 221.3 118.755 ;
      RECT 222.295 0.17 223.065 0.94 ;
      RECT 222.295 0.17 222.555 8.7 ;
      RECT 222.805 0.17 223.065 12.9 ;
      RECT 221.595 118.025 221.795 118.755 ;
      RECT 222.095 118.025 222.295 118.755 ;
      RECT 222.595 118.025 222.795 118.755 ;
      RECT 223.09 118.025 223.29 118.755 ;
      RECT 223.315 0.52 223.575 2.485 ;
      RECT 223.91 118.025 224.11 118.755 ;
      RECT 224.18 0.52 224.44 14.11 ;
      RECT 224.405 118.025 224.605 118.755 ;
      RECT 224.69 0.52 224.95 2.335 ;
      RECT 224.905 118.025 225.105 118.755 ;
      RECT 225.405 118.025 225.605 118.755 ;
      RECT 225.9 118.025 226.1 118.755 ;
      RECT 228.09 0.52 228.35 5.16 ;
      RECT 227.57 4.9 228.35 5.16 ;
      RECT 227.57 4.9 227.83 6.64 ;
      RECT 226.72 118.025 226.92 118.755 ;
      RECT 227.215 118.025 227.415 118.755 ;
      RECT 227.715 118.025 227.915 118.755 ;
      RECT 228.215 118.025 228.415 118.755 ;
      RECT 228.71 118.025 228.91 118.755 ;
      RECT 229.455 0.17 230.225 0.94 ;
      RECT 229.455 0.17 229.715 12.9 ;
      RECT 229.965 0.17 230.225 12.9 ;
      RECT 228.945 0.52 229.205 5.815 ;
      RECT 229.53 118.025 229.73 118.755 ;
      RECT 230.475 0.17 231.245 0.43 ;
      RECT 230.475 0.17 230.735 11.5 ;
      RECT 230.985 0.17 231.245 11.5 ;
      RECT 230.025 118.025 230.225 118.755 ;
      RECT 230.525 118.025 230.725 118.755 ;
      RECT 231.025 118.025 231.225 118.755 ;
      RECT 232.515 0.17 233.285 0.43 ;
      RECT 232.515 0.17 232.775 10.48 ;
      RECT 233.025 0.17 233.285 10.99 ;
      RECT 231.52 118.025 231.72 118.755 ;
      RECT 232.34 118.025 232.54 118.755 ;
      RECT 233.535 0.17 234.305 0.94 ;
      RECT 233.535 0.17 233.795 8.7 ;
      RECT 234.045 0.17 234.305 12.9 ;
      RECT 232.835 118.025 233.035 118.755 ;
      RECT 233.335 118.025 233.535 118.755 ;
      RECT 233.835 118.025 234.035 118.755 ;
      RECT 234.33 118.025 234.53 118.755 ;
      RECT 234.555 0.52 234.815 2.485 ;
      RECT 235.15 118.025 235.35 118.755 ;
      RECT 235.42 0.52 235.68 14.11 ;
      RECT 235.645 118.025 235.845 118.755 ;
      RECT 235.93 0.52 236.19 2.335 ;
      RECT 236.145 118.025 236.345 118.755 ;
      RECT 236.645 118.025 236.845 118.755 ;
      RECT 237.14 118.025 237.34 118.755 ;
      RECT 239.33 0.52 239.59 5.16 ;
      RECT 238.81 4.9 239.59 5.16 ;
      RECT 238.81 4.9 239.07 6.64 ;
      RECT 237.96 118.025 238.16 118.755 ;
      RECT 238.455 118.025 238.655 118.755 ;
      RECT 238.955 118.025 239.155 118.755 ;
      RECT 239.455 118.025 239.655 118.755 ;
      RECT 239.95 118.025 240.15 118.755 ;
      RECT 240.695 0.17 241.465 0.94 ;
      RECT 240.695 0.17 240.955 12.9 ;
      RECT 241.205 0.17 241.465 12.9 ;
      RECT 240.185 0.52 240.445 5.815 ;
      RECT 240.77 118.025 240.97 118.755 ;
      RECT 241.715 0.17 242.485 0.43 ;
      RECT 241.715 0.17 241.975 11.5 ;
      RECT 242.225 0.17 242.485 11.5 ;
      RECT 241.265 118.025 241.465 118.755 ;
      RECT 241.765 118.025 241.965 118.755 ;
      RECT 242.265 118.025 242.465 118.755 ;
      RECT 243.755 0.17 244.525 0.43 ;
      RECT 243.755 0.17 244.015 10.48 ;
      RECT 244.265 0.17 244.525 10.99 ;
      RECT 242.76 118.025 242.96 118.755 ;
      RECT 243.58 118.025 243.78 118.755 ;
      RECT 244.775 0.17 245.545 0.94 ;
      RECT 244.775 0.17 245.035 8.7 ;
      RECT 245.285 0.17 245.545 12.9 ;
      RECT 244.075 118.025 244.275 118.755 ;
      RECT 244.575 118.025 244.775 118.755 ;
      RECT 245.075 118.025 245.275 118.755 ;
      RECT 245.57 118.025 245.77 118.755 ;
      RECT 245.795 0.52 246.055 2.485 ;
      RECT 246.39 118.025 246.59 118.755 ;
      RECT 246.66 0.52 246.92 14.11 ;
      RECT 246.885 118.025 247.085 118.755 ;
      RECT 247.17 0.52 247.43 2.335 ;
      RECT 247.385 118.025 247.585 118.755 ;
      RECT 247.885 118.025 248.085 118.755 ;
      RECT 248.38 118.025 248.58 118.755 ;
      RECT 250.57 0.52 250.83 5.16 ;
      RECT 250.05 4.9 250.83 5.16 ;
      RECT 250.05 4.9 250.31 6.64 ;
      RECT 249.2 118.025 249.4 118.755 ;
      RECT 249.695 118.025 249.895 118.755 ;
      RECT 250.195 118.025 250.395 118.755 ;
      RECT 250.695 118.025 250.895 118.755 ;
      RECT 251.19 118.025 251.39 118.755 ;
      RECT 251.935 0.17 252.705 0.94 ;
      RECT 251.935 0.17 252.195 12.9 ;
      RECT 252.445 0.17 252.705 12.9 ;
      RECT 251.425 0.52 251.685 5.815 ;
      RECT 252.01 118.025 252.21 118.755 ;
      RECT 252.955 0.17 253.725 0.43 ;
      RECT 252.955 0.17 253.215 11.5 ;
      RECT 253.465 0.17 253.725 11.5 ;
      RECT 252.505 118.025 252.705 118.755 ;
      RECT 253.005 118.025 253.205 118.755 ;
      RECT 253.505 118.025 253.705 118.755 ;
      RECT 254.995 0.17 255.765 0.43 ;
      RECT 254.995 0.17 255.255 10.48 ;
      RECT 255.505 0.17 255.765 10.99 ;
      RECT 254 118.025 254.2 118.755 ;
      RECT 254.82 118.025 255.02 118.755 ;
      RECT 256.015 0.17 256.785 0.94 ;
      RECT 256.015 0.17 256.275 8.7 ;
      RECT 256.525 0.17 256.785 12.9 ;
      RECT 255.315 118.025 255.515 118.755 ;
      RECT 255.815 118.025 256.015 118.755 ;
      RECT 256.315 118.025 256.515 118.755 ;
      RECT 256.81 118.025 257.01 118.755 ;
      RECT 257.035 0.52 257.295 2.485 ;
      RECT 257.63 118.025 257.83 118.755 ;
      RECT 257.9 0.52 258.16 14.11 ;
      RECT 258.125 118.025 258.325 118.755 ;
      RECT 258.41 0.52 258.67 2.335 ;
      RECT 258.625 118.025 258.825 118.755 ;
      RECT 259.125 118.025 259.325 118.755 ;
      RECT 259.62 118.025 259.82 118.755 ;
      RECT 261.81 0.52 262.07 5.16 ;
      RECT 261.29 4.9 262.07 5.16 ;
      RECT 261.29 4.9 261.55 6.64 ;
      RECT 260.44 118.025 260.64 118.755 ;
      RECT 260.935 118.025 261.135 118.755 ;
      RECT 261.435 118.025 261.635 118.755 ;
      RECT 261.935 118.025 262.135 118.755 ;
      RECT 262.43 118.025 262.63 118.755 ;
      RECT 263.175 0.17 263.945 0.94 ;
      RECT 263.175 0.17 263.435 12.9 ;
      RECT 263.685 0.17 263.945 12.9 ;
      RECT 262.665 0.52 262.925 5.815 ;
      RECT 263.25 118.025 263.45 118.755 ;
      RECT 264.195 0.17 264.965 0.43 ;
      RECT 264.195 0.17 264.455 11.5 ;
      RECT 264.705 0.17 264.965 11.5 ;
      RECT 263.745 118.025 263.945 118.755 ;
      RECT 264.245 118.025 264.445 118.755 ;
      RECT 264.745 118.025 264.945 118.755 ;
      RECT 266.235 0.17 267.005 0.43 ;
      RECT 266.235 0.17 266.495 10.48 ;
      RECT 266.745 0.17 267.005 10.99 ;
      RECT 265.24 118.025 265.44 118.755 ;
      RECT 266.06 118.025 266.26 118.755 ;
      RECT 267.255 0.17 268.025 0.94 ;
      RECT 267.255 0.17 267.515 8.7 ;
      RECT 267.765 0.17 268.025 12.9 ;
      RECT 266.555 118.025 266.755 118.755 ;
      RECT 267.055 118.025 267.255 118.755 ;
      RECT 267.555 118.025 267.755 118.755 ;
      RECT 268.05 118.025 268.25 118.755 ;
      RECT 268.275 0.52 268.535 2.485 ;
      RECT 268.87 118.025 269.07 118.755 ;
      RECT 269.14 0.52 269.4 14.11 ;
      RECT 269.365 118.025 269.565 118.755 ;
      RECT 269.65 0.52 269.91 2.335 ;
      RECT 269.865 118.025 270.065 118.755 ;
      RECT 270.365 118.025 270.565 118.755 ;
      RECT 272.355 0.17 273.125 0.43 ;
      RECT 272.355 0.17 272.615 8.7 ;
      RECT 272.865 0.17 273.125 8.7 ;
      RECT 273.375 0.17 274.145 0.94 ;
      RECT 273.375 0.17 273.635 8.7 ;
      RECT 273.885 0.17 274.145 8.7 ;
      RECT 274.395 0.17 275.165 0.43 ;
      RECT 274.395 0.17 274.655 8.7 ;
      RECT 274.905 0.17 275.165 8.7 ;
      RECT 275.415 0.17 276.185 0.94 ;
      RECT 275.415 0.17 275.675 8.7 ;
      RECT 275.925 0.17 276.185 8.7 ;
      RECT 276.435 0.17 277.205 0.43 ;
      RECT 276.435 0.17 276.695 8.7 ;
      RECT 276.945 0.17 277.205 8.7 ;
      RECT 277.455 0.17 278.225 0.94 ;
      RECT 277.455 0.17 277.715 8.7 ;
      RECT 277.965 0.17 278.225 8.7 ;
      RECT 270.86 118.025 271.06 118.755 ;
      RECT 271.68 118.025 271.88 118.755 ;
      RECT 272.675 118.025 272.875 118.755 ;
      RECT 280.16 0.17 280.93 0.94 ;
      RECT 280.16 0.17 280.42 8.7 ;
      RECT 280.67 0.17 280.93 8.7 ;
      RECT 278.63 0.3 278.89 8.7 ;
      RECT 279.14 0 279.4 8.7 ;
      RECT 279.65 0 279.91 8.7 ;
      RECT 281.18 0 281.44 8.7 ;
      RECT 281.69 0 281.95 8.7 ;
      RECT 282.2 0.52 282.46 8.7 ;
      RECT 282.71 0.52 282.97 8.7 ;
      RECT 283.22 0.52 283.48 8.7 ;
      RECT 285.26 0.17 286.03 0.94 ;
      RECT 285.26 0.17 285.52 8.7 ;
      RECT 285.77 0.17 286.03 8.7 ;
      RECT 286.28 0.17 287.05 0.43 ;
      RECT 286.28 0.17 286.54 8.7 ;
      RECT 286.79 0.17 287.05 8.7 ;
      RECT 283.73 0.52 283.99 8.7 ;
      RECT 284.24 0 284.5 8.7 ;
      RECT 284.75 0 285.01 8.7 ;
      RECT 287.3 0.3 287.56 8.7 ;
      RECT 287.81 0.3 288.07 8.7 ;
      RECT 289.85 0.17 290.62 0.94 ;
      RECT 289.85 0.17 290.11 8.7 ;
      RECT 290.36 0.17 290.62 8.7 ;
      RECT 288.32 0.3 288.58 8.7 ;
      RECT 288.83 0.3 289.09 8.7 ;
      RECT 289.34 0.3 289.6 8.7 ;
      RECT 290.87 0.52 291.13 8.7 ;
      RECT 291.38 0.52 291.64 8.7 ;
      RECT 291.89 0.3 292.15 8.7 ;
      RECT 292.4 0.52 292.66 8.7 ;
      RECT 292.91 0.52 293.17 8.7 ;
      RECT 293.42 0.3 293.68 8.7 ;
      RECT 293.93 0.52 294.19 8.7 ;
      RECT 294.44 0.52 294.7 8.7 ;
      RECT 294.95 0.52 295.21 8.7 ;
      RECT 295.46 0.52 295.72 8.7 ;
      RECT 295.97 0.52 296.23 8.7 ;
      RECT 296.48 0.3 296.74 8.7 ;
      RECT 296.99 0.52 297.25 8.7 ;
      RECT 297.5 0.52 297.76 8.7 ;
      RECT 298.01 0.3 298.27 8.7 ;
      RECT 300.05 0.17 300.82 0.94 ;
      RECT 300.05 0.17 300.31 8.7 ;
      RECT 300.56 0.17 300.82 8.7 ;
      RECT 298.52 0.52 298.78 8.7 ;
      RECT 299.03 0.52 299.29 8.7 ;
      RECT 299.54 0.3 299.8 8.7 ;
      RECT 301.07 0.52 301.33 8.7 ;
      RECT 301.58 0.52 301.84 8.7 ;
      RECT 302.09 0.52 302.35 8.7 ;
      RECT 302.6 0.52 302.86 8.7 ;
      RECT 303.11 0.52 303.37 8.7 ;
      RECT 303.62 0.52 303.88 8.7 ;
      RECT 304.13 0.52 304.39 8.7 ;
      RECT 306.17 0.17 306.94 0.94 ;
      RECT 306.17 0.17 306.43 8.7 ;
      RECT 306.68 0.17 306.94 8.7 ;
      RECT 304.64 0.52 304.9 8.7 ;
      RECT 305.15 0 305.41 8.7 ;
      RECT 305.66 0 305.92 8.7 ;
      RECT 307.19 0 307.45 8.7 ;
      RECT 309.23 0.17 310 0.43 ;
      RECT 309.23 0.17 309.49 8.7 ;
      RECT 309.74 0.17 310 8.7 ;
      RECT 307.7 0 307.96 8.7 ;
      RECT 308.21 0.3 308.47 8.7 ;
      RECT 308.72 0.3 308.98 8.7 ;
      RECT 310.25 0.3 310.51 8.7 ;
      RECT 310.76 0.3 311.02 8.7 ;
      RECT 311.27 0.3 311.53 8.7 ;
      RECT 311.78 0.3 312.04 8.7 ;
      RECT 312.29 0 312.55 8.7 ;
      RECT 312.8 0 313.06 8.7 ;
      RECT 314.84 0.17 315.61 0.43 ;
      RECT 314.84 0.17 315.1 8.7 ;
      RECT 315.35 0.17 315.61 8.7 ;
      RECT 315.86 0.17 316.63 0.94 ;
      RECT 315.86 0.17 316.12 25.5 ;
      RECT 316.37 0.17 316.63 33.9 ;
      RECT 316.88 0.17 317.65 0.43 ;
      RECT 316.88 0.17 317.14 8.7 ;
      RECT 317.39 0.17 317.65 8.7 ;
      RECT 318.255 0.17 319.025 0.94 ;
      RECT 318.255 0.17 318.515 8.7 ;
      RECT 318.765 0.17 319.025 8.7 ;
      RECT 319.275 0.17 320.045 0.43 ;
      RECT 319.275 0.17 319.535 8.7 ;
      RECT 319.785 0.17 320.045 8.7 ;
      RECT 320.295 0.17 321.065 0.94 ;
      RECT 320.295 0.17 320.555 8.7 ;
      RECT 320.805 0.17 321.065 8.7 ;
      RECT 321.315 0.17 322.085 0.43 ;
      RECT 321.315 0.17 321.575 8.7 ;
      RECT 321.825 0.17 322.085 8.7 ;
      RECT 322.335 0.17 323.105 0.94 ;
      RECT 322.335 0.17 322.595 8.7 ;
      RECT 322.845 0.17 323.105 8.7 ;
      RECT 313.31 0.3 313.57 8.7 ;
      RECT 323.355 0.17 324.125 0.43 ;
      RECT 323.355 0.17 323.615 8.7 ;
      RECT 323.865 0.17 324.125 8.7 ;
      RECT 313.82 0.3 314.08 8.7 ;
      RECT 314.33 0.52 314.59 8.7 ;
      RECT 323.605 118.025 323.805 118.755 ;
      RECT 324.6 118.025 324.8 118.755 ;
      RECT 325.42 118.025 325.62 118.755 ;
      RECT 325.915 118.025 326.115 118.755 ;
      RECT 326.415 118.025 326.615 118.755 ;
      RECT 326.57 0.52 326.83 2.335 ;
      RECT 326.915 118.025 327.115 118.755 ;
      RECT 327.08 0.52 327.34 14.11 ;
      RECT 327.41 118.025 327.61 118.755 ;
      RECT 328.455 0.17 329.225 0.94 ;
      RECT 328.965 0.17 329.225 8.7 ;
      RECT 328.455 0.17 328.715 12.9 ;
      RECT 327.945 0.52 328.205 2.485 ;
      RECT 328.23 118.025 328.43 118.755 ;
      RECT 329.475 0.17 330.245 0.43 ;
      RECT 329.985 0.17 330.245 10.48 ;
      RECT 329.475 0.17 329.735 10.99 ;
      RECT 328.725 118.025 328.925 118.755 ;
      RECT 329.225 118.025 329.425 118.755 ;
      RECT 329.725 118.025 329.925 118.755 ;
      RECT 330.22 118.025 330.42 118.755 ;
      RECT 331.515 0.17 332.285 0.43 ;
      RECT 331.515 0.17 331.775 11.5 ;
      RECT 332.025 0.17 332.285 11.5 ;
      RECT 331.04 118.025 331.24 118.755 ;
      RECT 331.535 118.025 331.735 118.755 ;
      RECT 332.535 0.17 333.305 0.94 ;
      RECT 332.535 0.17 332.795 12.9 ;
      RECT 333.045 0.17 333.305 12.9 ;
      RECT 332.035 118.025 332.235 118.755 ;
      RECT 332.535 118.025 332.735 118.755 ;
      RECT 333.03 118.025 333.23 118.755 ;
      RECT 333.555 0.52 333.815 5.815 ;
      RECT 334.41 0.52 334.67 5.16 ;
      RECT 334.41 4.9 335.19 5.16 ;
      RECT 334.93 4.9 335.19 6.64 ;
      RECT 333.85 118.025 334.05 118.755 ;
      RECT 334.345 118.025 334.545 118.755 ;
      RECT 334.845 118.025 335.045 118.755 ;
      RECT 335.345 118.025 335.545 118.755 ;
      RECT 335.84 118.025 336.04 118.755 ;
      RECT 336.66 118.025 336.86 118.755 ;
      RECT 337.155 118.025 337.355 118.755 ;
      RECT 337.655 118.025 337.855 118.755 ;
      RECT 337.81 0.52 338.07 2.335 ;
      RECT 338.155 118.025 338.355 118.755 ;
      RECT 338.32 0.52 338.58 14.11 ;
      RECT 338.65 118.025 338.85 118.755 ;
      RECT 339.695 0.17 340.465 0.94 ;
      RECT 340.205 0.17 340.465 8.7 ;
      RECT 339.695 0.17 339.955 12.9 ;
      RECT 339.185 0.52 339.445 2.485 ;
      RECT 339.47 118.025 339.67 118.755 ;
      RECT 340.715 0.17 341.485 0.43 ;
      RECT 341.225 0.17 341.485 10.48 ;
      RECT 340.715 0.17 340.975 10.99 ;
      RECT 339.965 118.025 340.165 118.755 ;
      RECT 340.465 118.025 340.665 118.755 ;
      RECT 340.965 118.025 341.165 118.755 ;
      RECT 341.46 118.025 341.66 118.755 ;
      RECT 342.755 0.17 343.525 0.43 ;
      RECT 342.755 0.17 343.015 11.5 ;
      RECT 343.265 0.17 343.525 11.5 ;
      RECT 342.28 118.025 342.48 118.755 ;
      RECT 342.775 118.025 342.975 118.755 ;
      RECT 343.775 0.17 344.545 0.94 ;
      RECT 343.775 0.17 344.035 12.9 ;
      RECT 344.285 0.17 344.545 12.9 ;
      RECT 343.275 118.025 343.475 118.755 ;
      RECT 343.775 118.025 343.975 118.755 ;
      RECT 344.27 118.025 344.47 118.755 ;
      RECT 344.795 0.52 345.055 5.815 ;
      RECT 345.65 0.52 345.91 5.16 ;
      RECT 345.65 4.9 346.43 5.16 ;
      RECT 346.17 4.9 346.43 6.64 ;
      RECT 345.09 118.025 345.29 118.755 ;
      RECT 345.585 118.025 345.785 118.755 ;
      RECT 346.085 118.025 346.285 118.755 ;
      RECT 346.585 118.025 346.785 118.755 ;
      RECT 347.08 118.025 347.28 118.755 ;
      RECT 347.9 118.025 348.1 118.755 ;
      RECT 348.395 118.025 348.595 118.755 ;
      RECT 348.895 118.025 349.095 118.755 ;
      RECT 349.05 0.52 349.31 2.335 ;
      RECT 349.395 118.025 349.595 118.755 ;
      RECT 349.56 0.52 349.82 14.11 ;
      RECT 349.89 118.025 350.09 118.755 ;
      RECT 350.935 0.17 351.705 0.94 ;
      RECT 351.445 0.17 351.705 8.7 ;
      RECT 350.935 0.17 351.195 12.9 ;
      RECT 350.425 0.52 350.685 2.485 ;
      RECT 350.71 118.025 350.91 118.755 ;
      RECT 351.955 0.17 352.725 0.43 ;
      RECT 352.465 0.17 352.725 10.48 ;
      RECT 351.955 0.17 352.215 10.99 ;
      RECT 351.205 118.025 351.405 118.755 ;
      RECT 351.705 118.025 351.905 118.755 ;
      RECT 352.205 118.025 352.405 118.755 ;
      RECT 352.7 118.025 352.9 118.755 ;
      RECT 353.995 0.17 354.765 0.43 ;
      RECT 353.995 0.17 354.255 11.5 ;
      RECT 354.505 0.17 354.765 11.5 ;
      RECT 353.52 118.025 353.72 118.755 ;
      RECT 354.015 118.025 354.215 118.755 ;
      RECT 355.015 0.17 355.785 0.94 ;
      RECT 355.015 0.17 355.275 12.9 ;
      RECT 355.525 0.17 355.785 12.9 ;
      RECT 354.515 118.025 354.715 118.755 ;
      RECT 355.015 118.025 355.215 118.755 ;
      RECT 355.51 118.025 355.71 118.755 ;
      RECT 356.035 0.52 356.295 5.815 ;
      RECT 356.89 0.52 357.15 5.16 ;
      RECT 356.89 4.9 357.67 5.16 ;
      RECT 357.41 4.9 357.67 6.64 ;
      RECT 356.33 118.025 356.53 118.755 ;
      RECT 356.825 118.025 357.025 118.755 ;
      RECT 357.325 118.025 357.525 118.755 ;
      RECT 357.825 118.025 358.025 118.755 ;
      RECT 358.32 118.025 358.52 118.755 ;
      RECT 359.14 118.025 359.34 118.755 ;
      RECT 359.635 118.025 359.835 118.755 ;
      RECT 360.135 118.025 360.335 118.755 ;
      RECT 360.29 0.52 360.55 2.335 ;
      RECT 360.635 118.025 360.835 118.755 ;
      RECT 360.8 0.52 361.06 14.11 ;
      RECT 361.13 118.025 361.33 118.755 ;
      RECT 362.175 0.17 362.945 0.94 ;
      RECT 362.685 0.17 362.945 8.7 ;
      RECT 362.175 0.17 362.435 12.9 ;
      RECT 361.665 0.52 361.925 2.485 ;
      RECT 361.95 118.025 362.15 118.755 ;
      RECT 363.195 0.17 363.965 0.43 ;
      RECT 363.705 0.17 363.965 10.48 ;
      RECT 363.195 0.17 363.455 10.99 ;
      RECT 362.445 118.025 362.645 118.755 ;
      RECT 362.945 118.025 363.145 118.755 ;
      RECT 363.445 118.025 363.645 118.755 ;
      RECT 363.94 118.025 364.14 118.755 ;
      RECT 365.235 0.17 366.005 0.43 ;
      RECT 365.235 0.17 365.495 11.5 ;
      RECT 365.745 0.17 366.005 11.5 ;
      RECT 364.76 118.025 364.96 118.755 ;
      RECT 365.255 118.025 365.455 118.755 ;
      RECT 366.255 0.17 367.025 0.94 ;
      RECT 366.255 0.17 366.515 12.9 ;
      RECT 366.765 0.17 367.025 12.9 ;
      RECT 365.755 118.025 365.955 118.755 ;
      RECT 366.255 118.025 366.455 118.755 ;
      RECT 366.75 118.025 366.95 118.755 ;
      RECT 367.275 0.52 367.535 5.815 ;
      RECT 368.13 0.52 368.39 5.16 ;
      RECT 368.13 4.9 368.91 5.16 ;
      RECT 368.65 4.9 368.91 6.64 ;
      RECT 367.57 118.025 367.77 118.755 ;
      RECT 368.065 118.025 368.265 118.755 ;
      RECT 368.565 118.025 368.765 118.755 ;
      RECT 369.065 118.025 369.265 118.755 ;
      RECT 369.56 118.025 369.76 118.755 ;
      RECT 370.38 118.025 370.58 118.755 ;
      RECT 370.875 118.025 371.075 118.755 ;
      RECT 371.375 118.025 371.575 118.755 ;
      RECT 371.53 0.52 371.79 2.335 ;
      RECT 371.875 118.025 372.075 118.755 ;
      RECT 372.04 0.52 372.3 14.11 ;
      RECT 372.37 118.025 372.57 118.755 ;
      RECT 373.415 0.17 374.185 0.94 ;
      RECT 373.925 0.17 374.185 8.7 ;
      RECT 373.415 0.17 373.675 12.9 ;
      RECT 372.905 0.52 373.165 2.485 ;
      RECT 373.19 118.025 373.39 118.755 ;
      RECT 374.435 0.17 375.205 0.43 ;
      RECT 374.945 0.17 375.205 10.48 ;
      RECT 374.435 0.17 374.695 10.99 ;
      RECT 373.685 118.025 373.885 118.755 ;
      RECT 374.185 118.025 374.385 118.755 ;
      RECT 374.685 118.025 374.885 118.755 ;
      RECT 375.18 118.025 375.38 118.755 ;
      RECT 376.475 0.17 377.245 0.43 ;
      RECT 376.475 0.17 376.735 11.5 ;
      RECT 376.985 0.17 377.245 11.5 ;
      RECT 376 118.025 376.2 118.755 ;
      RECT 376.495 118.025 376.695 118.755 ;
      RECT 377.495 0.17 378.265 0.94 ;
      RECT 377.495 0.17 377.755 12.9 ;
      RECT 378.005 0.17 378.265 12.9 ;
      RECT 376.995 118.025 377.195 118.755 ;
      RECT 377.495 118.025 377.695 118.755 ;
      RECT 377.99 118.025 378.19 118.755 ;
      RECT 378.515 0.52 378.775 5.815 ;
      RECT 379.37 0.52 379.63 5.16 ;
      RECT 379.37 4.9 380.15 5.16 ;
      RECT 379.89 4.9 380.15 6.64 ;
      RECT 378.81 118.025 379.01 118.755 ;
      RECT 379.305 118.025 379.505 118.755 ;
      RECT 379.805 118.025 380.005 118.755 ;
      RECT 380.305 118.025 380.505 118.755 ;
      RECT 380.8 118.025 381 118.755 ;
      RECT 381.62 118.025 381.82 118.755 ;
      RECT 382.115 118.025 382.315 118.755 ;
      RECT 382.615 118.025 382.815 118.755 ;
      RECT 382.77 0.52 383.03 2.335 ;
      RECT 383.115 118.025 383.315 118.755 ;
      RECT 383.28 0.52 383.54 14.11 ;
      RECT 383.61 118.025 383.81 118.755 ;
      RECT 384.655 0.17 385.425 0.94 ;
      RECT 385.165 0.17 385.425 8.7 ;
      RECT 384.655 0.17 384.915 12.9 ;
      RECT 384.145 0.52 384.405 2.485 ;
      RECT 384.43 118.025 384.63 118.755 ;
      RECT 385.675 0.17 386.445 0.43 ;
      RECT 386.185 0.17 386.445 10.48 ;
      RECT 385.675 0.17 385.935 10.99 ;
      RECT 384.925 118.025 385.125 118.755 ;
      RECT 385.425 118.025 385.625 118.755 ;
      RECT 385.925 118.025 386.125 118.755 ;
      RECT 386.42 118.025 386.62 118.755 ;
      RECT 387.715 0.17 388.485 0.43 ;
      RECT 387.715 0.17 387.975 11.5 ;
      RECT 388.225 0.17 388.485 11.5 ;
      RECT 387.24 118.025 387.44 118.755 ;
      RECT 387.735 118.025 387.935 118.755 ;
      RECT 388.735 0.17 389.505 0.94 ;
      RECT 388.735 0.17 388.995 12.9 ;
      RECT 389.245 0.17 389.505 12.9 ;
      RECT 388.235 118.025 388.435 118.755 ;
      RECT 388.735 118.025 388.935 118.755 ;
      RECT 389.23 118.025 389.43 118.755 ;
      RECT 389.755 0.52 390.015 5.815 ;
      RECT 390.61 0.52 390.87 5.16 ;
      RECT 390.61 4.9 391.39 5.16 ;
      RECT 391.13 4.9 391.39 6.64 ;
      RECT 390.05 118.025 390.25 118.755 ;
      RECT 390.545 118.025 390.745 118.755 ;
      RECT 391.045 118.025 391.245 118.755 ;
      RECT 391.545 118.025 391.745 118.755 ;
      RECT 392.04 118.025 392.24 118.755 ;
      RECT 392.86 118.025 393.06 118.755 ;
      RECT 393.355 118.025 393.555 118.755 ;
      RECT 393.855 118.025 394.055 118.755 ;
      RECT 394.01 0.52 394.27 2.335 ;
      RECT 394.355 118.025 394.555 118.755 ;
      RECT 394.52 0.52 394.78 14.11 ;
      RECT 394.85 118.025 395.05 118.755 ;
      RECT 395.895 0.17 396.665 0.94 ;
      RECT 396.405 0.17 396.665 8.7 ;
      RECT 395.895 0.17 396.155 12.9 ;
      RECT 395.385 0.52 395.645 2.485 ;
      RECT 395.67 118.025 395.87 118.755 ;
      RECT 396.915 0.17 397.685 0.43 ;
      RECT 397.425 0.17 397.685 10.48 ;
      RECT 396.915 0.17 397.175 10.99 ;
      RECT 396.165 118.025 396.365 118.755 ;
      RECT 396.665 118.025 396.865 118.755 ;
      RECT 397.165 118.025 397.365 118.755 ;
      RECT 397.66 118.025 397.86 118.755 ;
      RECT 398.955 0.17 399.725 0.43 ;
      RECT 398.955 0.17 399.215 11.5 ;
      RECT 399.465 0.17 399.725 11.5 ;
      RECT 398.48 118.025 398.68 118.755 ;
      RECT 398.975 118.025 399.175 118.755 ;
      RECT 399.975 0.17 400.745 0.94 ;
      RECT 399.975 0.17 400.235 12.9 ;
      RECT 400.485 0.17 400.745 12.9 ;
      RECT 399.475 118.025 399.675 118.755 ;
      RECT 399.975 118.025 400.175 118.755 ;
      RECT 400.47 118.025 400.67 118.755 ;
      RECT 400.995 0.52 401.255 5.815 ;
      RECT 401.85 0.52 402.11 5.16 ;
      RECT 401.85 4.9 402.63 5.16 ;
      RECT 402.37 4.9 402.63 6.64 ;
      RECT 401.29 118.025 401.49 118.755 ;
      RECT 401.785 118.025 401.985 118.755 ;
      RECT 402.285 118.025 402.485 118.755 ;
      RECT 402.785 118.025 402.985 118.755 ;
      RECT 403.28 118.025 403.48 118.755 ;
      RECT 404.1 118.025 404.3 118.755 ;
      RECT 404.595 118.025 404.795 118.755 ;
      RECT 405.095 118.025 405.295 118.755 ;
      RECT 405.25 0.52 405.51 2.335 ;
      RECT 405.595 118.025 405.795 118.755 ;
      RECT 405.76 0.52 406.02 14.11 ;
      RECT 406.09 118.025 406.29 118.755 ;
      RECT 407.135 0.17 407.905 0.94 ;
      RECT 407.645 0.17 407.905 8.7 ;
      RECT 407.135 0.17 407.395 12.9 ;
      RECT 406.625 0.52 406.885 2.485 ;
      RECT 406.91 118.025 407.11 118.755 ;
      RECT 408.155 0.17 408.925 0.43 ;
      RECT 408.665 0.17 408.925 10.48 ;
      RECT 408.155 0.17 408.415 10.99 ;
      RECT 407.405 118.025 407.605 118.755 ;
      RECT 407.905 118.025 408.105 118.755 ;
      RECT 408.405 118.025 408.605 118.755 ;
      RECT 408.9 118.025 409.1 118.755 ;
      RECT 410.195 0.17 410.965 0.43 ;
      RECT 410.195 0.17 410.455 11.5 ;
      RECT 410.705 0.17 410.965 11.5 ;
      RECT 409.72 118.025 409.92 118.755 ;
      RECT 410.215 118.025 410.415 118.755 ;
      RECT 411.215 0.17 411.985 0.94 ;
      RECT 411.215 0.17 411.475 12.9 ;
      RECT 411.725 0.17 411.985 12.9 ;
      RECT 410.715 118.025 410.915 118.755 ;
      RECT 411.215 118.025 411.415 118.755 ;
      RECT 411.71 118.025 411.91 118.755 ;
      RECT 412.235 0.52 412.495 5.815 ;
      RECT 413.09 0.52 413.35 5.16 ;
      RECT 413.09 4.9 413.87 5.16 ;
      RECT 413.61 4.9 413.87 6.64 ;
      RECT 412.53 118.025 412.73 118.755 ;
      RECT 413.025 118.025 413.225 118.755 ;
      RECT 413.525 118.025 413.725 118.755 ;
      RECT 414.025 118.025 414.225 118.755 ;
      RECT 414.52 118.025 414.72 118.755 ;
      RECT 415.34 118.025 415.54 118.755 ;
      RECT 415.835 118.025 416.035 118.755 ;
      RECT 416.335 118.025 416.535 118.755 ;
      RECT 416.49 0.52 416.75 2.335 ;
      RECT 416.835 118.025 417.035 118.755 ;
      RECT 417 0.52 417.26 14.11 ;
      RECT 417.33 118.025 417.53 118.755 ;
      RECT 418.375 0.17 419.145 0.94 ;
      RECT 418.885 0.17 419.145 8.7 ;
      RECT 418.375 0.17 418.635 12.9 ;
      RECT 417.865 0.52 418.125 2.485 ;
      RECT 418.15 118.025 418.35 118.755 ;
      RECT 419.395 0.17 420.165 0.43 ;
      RECT 419.905 0.17 420.165 10.48 ;
      RECT 419.395 0.17 419.655 10.99 ;
      RECT 418.645 118.025 418.845 118.755 ;
      RECT 419.145 118.025 419.345 118.755 ;
      RECT 419.645 118.025 419.845 118.755 ;
      RECT 420.14 118.025 420.34 118.755 ;
      RECT 421.435 0.17 422.205 0.43 ;
      RECT 421.435 0.17 421.695 11.5 ;
      RECT 421.945 0.17 422.205 11.5 ;
      RECT 420.96 118.025 421.16 118.755 ;
      RECT 421.455 118.025 421.655 118.755 ;
      RECT 422.455 0.17 423.225 0.94 ;
      RECT 422.455 0.17 422.715 12.9 ;
      RECT 422.965 0.17 423.225 12.9 ;
      RECT 421.955 118.025 422.155 118.755 ;
      RECT 422.455 118.025 422.655 118.755 ;
      RECT 422.95 118.025 423.15 118.755 ;
      RECT 423.475 0.52 423.735 5.815 ;
      RECT 424.33 0.52 424.59 5.16 ;
      RECT 424.33 4.9 425.11 5.16 ;
      RECT 424.85 4.9 425.11 6.64 ;
      RECT 423.77 118.025 423.97 118.755 ;
      RECT 424.265 118.025 424.465 118.755 ;
      RECT 424.765 118.025 424.965 118.755 ;
      RECT 425.265 118.025 425.465 118.755 ;
      RECT 425.76 118.025 425.96 118.755 ;
      RECT 426.58 118.025 426.78 118.755 ;
      RECT 427.075 118.025 427.275 118.755 ;
      RECT 427.575 118.025 427.775 118.755 ;
      RECT 427.73 0.52 427.99 2.335 ;
      RECT 428.075 118.025 428.275 118.755 ;
      RECT 428.24 0.52 428.5 14.11 ;
      RECT 428.57 118.025 428.77 118.755 ;
      RECT 429.615 0.17 430.385 0.94 ;
      RECT 430.125 0.17 430.385 8.7 ;
      RECT 429.615 0.17 429.875 12.9 ;
      RECT 429.105 0.52 429.365 2.485 ;
      RECT 429.39 118.025 429.59 118.755 ;
      RECT 430.635 0.17 431.405 0.43 ;
      RECT 431.145 0.17 431.405 10.48 ;
      RECT 430.635 0.17 430.895 10.99 ;
      RECT 429.885 118.025 430.085 118.755 ;
      RECT 430.385 118.025 430.585 118.755 ;
      RECT 430.885 118.025 431.085 118.755 ;
      RECT 431.38 118.025 431.58 118.755 ;
      RECT 432.675 0.17 433.445 0.43 ;
      RECT 432.675 0.17 432.935 11.5 ;
      RECT 433.185 0.17 433.445 11.5 ;
      RECT 432.2 118.025 432.4 118.755 ;
      RECT 432.695 118.025 432.895 118.755 ;
      RECT 433.695 0.17 434.465 0.94 ;
      RECT 433.695 0.17 433.955 12.9 ;
      RECT 434.205 0.17 434.465 12.9 ;
      RECT 433.195 118.025 433.395 118.755 ;
      RECT 433.695 118.025 433.895 118.755 ;
      RECT 434.19 118.025 434.39 118.755 ;
      RECT 434.715 0.52 434.975 5.815 ;
      RECT 435.57 0.52 435.83 5.16 ;
      RECT 435.57 4.9 436.35 5.16 ;
      RECT 436.09 4.9 436.35 6.64 ;
      RECT 435.01 118.025 435.21 118.755 ;
      RECT 435.505 118.025 435.705 118.755 ;
      RECT 436.005 118.025 436.205 118.755 ;
      RECT 436.505 118.025 436.705 118.755 ;
      RECT 437 118.025 437.2 118.755 ;
      RECT 437.82 118.025 438.02 118.755 ;
      RECT 438.315 118.025 438.515 118.755 ;
      RECT 438.815 118.025 439.015 118.755 ;
      RECT 438.97 0.52 439.23 2.335 ;
      RECT 439.315 118.025 439.515 118.755 ;
      RECT 439.48 0.52 439.74 14.11 ;
      RECT 439.81 118.025 440.01 118.755 ;
      RECT 440.855 0.17 441.625 0.94 ;
      RECT 441.365 0.17 441.625 8.7 ;
      RECT 440.855 0.17 441.115 12.9 ;
      RECT 440.345 0.52 440.605 2.485 ;
      RECT 440.63 118.025 440.83 118.755 ;
      RECT 441.875 0.17 442.645 0.43 ;
      RECT 442.385 0.17 442.645 10.48 ;
      RECT 441.875 0.17 442.135 10.99 ;
      RECT 441.125 118.025 441.325 118.755 ;
      RECT 441.625 118.025 441.825 118.755 ;
      RECT 442.125 118.025 442.325 118.755 ;
      RECT 442.62 118.025 442.82 118.755 ;
      RECT 443.915 0.17 444.685 0.43 ;
      RECT 443.915 0.17 444.175 11.5 ;
      RECT 444.425 0.17 444.685 11.5 ;
      RECT 443.44 118.025 443.64 118.755 ;
      RECT 443.935 118.025 444.135 118.755 ;
      RECT 444.935 0.17 445.705 0.94 ;
      RECT 444.935 0.17 445.195 12.9 ;
      RECT 445.445 0.17 445.705 12.9 ;
      RECT 444.435 118.025 444.635 118.755 ;
      RECT 444.935 118.025 445.135 118.755 ;
      RECT 445.43 118.025 445.63 118.755 ;
      RECT 445.955 0.52 446.215 5.815 ;
      RECT 446.81 0.52 447.07 5.16 ;
      RECT 446.81 4.9 447.59 5.16 ;
      RECT 447.33 4.9 447.59 6.64 ;
      RECT 446.25 118.025 446.45 118.755 ;
      RECT 446.745 118.025 446.945 118.755 ;
      RECT 447.245 118.025 447.445 118.755 ;
      RECT 447.745 118.025 447.945 118.755 ;
      RECT 448.24 118.025 448.44 118.755 ;
      RECT 449.06 118.025 449.26 118.755 ;
      RECT 449.555 118.025 449.755 118.755 ;
      RECT 450.055 118.025 450.255 118.755 ;
      RECT 450.21 0.52 450.47 2.335 ;
      RECT 450.555 118.025 450.755 118.755 ;
      RECT 450.72 0.52 450.98 14.11 ;
      RECT 451.05 118.025 451.25 118.755 ;
      RECT 452.095 0.17 452.865 0.94 ;
      RECT 452.605 0.17 452.865 8.7 ;
      RECT 452.095 0.17 452.355 12.9 ;
      RECT 451.585 0.52 451.845 2.485 ;
      RECT 451.87 118.025 452.07 118.755 ;
      RECT 453.115 0.17 453.885 0.43 ;
      RECT 453.625 0.17 453.885 10.48 ;
      RECT 453.115 0.17 453.375 10.99 ;
      RECT 452.365 118.025 452.565 118.755 ;
      RECT 452.865 118.025 453.065 118.755 ;
      RECT 453.365 118.025 453.565 118.755 ;
      RECT 453.86 118.025 454.06 118.755 ;
      RECT 455.155 0.17 455.925 0.43 ;
      RECT 455.155 0.17 455.415 11.5 ;
      RECT 455.665 0.17 455.925 11.5 ;
      RECT 454.68 118.025 454.88 118.755 ;
      RECT 455.175 118.025 455.375 118.755 ;
      RECT 456.175 0.17 456.945 0.94 ;
      RECT 456.175 0.17 456.435 12.9 ;
      RECT 456.685 0.17 456.945 12.9 ;
      RECT 455.675 118.025 455.875 118.755 ;
      RECT 456.175 118.025 456.375 118.755 ;
      RECT 456.67 118.025 456.87 118.755 ;
      RECT 457.195 0.52 457.455 5.815 ;
      RECT 458.05 0.52 458.31 5.16 ;
      RECT 458.05 4.9 458.83 5.16 ;
      RECT 458.57 4.9 458.83 6.64 ;
      RECT 457.49 118.025 457.69 118.755 ;
      RECT 457.985 118.025 458.185 118.755 ;
      RECT 458.485 118.025 458.685 118.755 ;
      RECT 458.985 118.025 459.185 118.755 ;
      RECT 459.48 118.025 459.68 118.755 ;
      RECT 460.3 118.025 460.5 118.755 ;
      RECT 460.795 118.025 460.995 118.755 ;
      RECT 461.295 118.025 461.495 118.755 ;
      RECT 461.45 0.52 461.71 2.335 ;
      RECT 461.795 118.025 461.995 118.755 ;
      RECT 461.96 0.52 462.22 14.11 ;
      RECT 462.29 118.025 462.49 118.755 ;
      RECT 463.335 0.17 464.105 0.94 ;
      RECT 463.845 0.17 464.105 8.7 ;
      RECT 463.335 0.17 463.595 12.9 ;
      RECT 462.825 0.52 463.085 2.485 ;
      RECT 463.11 118.025 463.31 118.755 ;
      RECT 464.355 0.17 465.125 0.43 ;
      RECT 464.865 0.17 465.125 10.48 ;
      RECT 464.355 0.17 464.615 10.99 ;
      RECT 463.605 118.025 463.805 118.755 ;
      RECT 464.105 118.025 464.305 118.755 ;
      RECT 464.605 118.025 464.805 118.755 ;
      RECT 465.1 118.025 465.3 118.755 ;
      RECT 466.395 0.17 467.165 0.43 ;
      RECT 466.395 0.17 466.655 11.5 ;
      RECT 466.905 0.17 467.165 11.5 ;
      RECT 465.92 118.025 466.12 118.755 ;
      RECT 466.415 118.025 466.615 118.755 ;
      RECT 467.415 0.17 468.185 0.94 ;
      RECT 467.415 0.17 467.675 12.9 ;
      RECT 467.925 0.17 468.185 12.9 ;
      RECT 466.915 118.025 467.115 118.755 ;
      RECT 467.415 118.025 467.615 118.755 ;
      RECT 467.91 118.025 468.11 118.755 ;
      RECT 468.435 0.52 468.695 5.815 ;
      RECT 469.29 0.52 469.55 5.16 ;
      RECT 469.29 4.9 470.07 5.16 ;
      RECT 469.81 4.9 470.07 6.64 ;
      RECT 468.73 118.025 468.93 118.755 ;
      RECT 469.225 118.025 469.425 118.755 ;
      RECT 469.725 118.025 469.925 118.755 ;
      RECT 470.225 118.025 470.425 118.755 ;
      RECT 470.72 118.025 470.92 118.755 ;
      RECT 471.54 118.025 471.74 118.755 ;
      RECT 472.035 118.025 472.235 118.755 ;
      RECT 472.535 118.025 472.735 118.755 ;
      RECT 472.69 0.52 472.95 2.335 ;
      RECT 473.035 118.025 473.235 118.755 ;
      RECT 473.2 0.52 473.46 14.11 ;
      RECT 473.53 118.025 473.73 118.755 ;
      RECT 474.575 0.17 475.345 0.94 ;
      RECT 475.085 0.17 475.345 8.7 ;
      RECT 474.575 0.17 474.835 12.9 ;
      RECT 474.065 0.52 474.325 2.485 ;
      RECT 474.35 118.025 474.55 118.755 ;
      RECT 475.595 0.17 476.365 0.43 ;
      RECT 476.105 0.17 476.365 10.48 ;
      RECT 475.595 0.17 475.855 10.99 ;
      RECT 474.845 118.025 475.045 118.755 ;
      RECT 475.345 118.025 475.545 118.755 ;
      RECT 475.845 118.025 476.045 118.755 ;
      RECT 476.34 118.025 476.54 118.755 ;
      RECT 477.635 0.17 478.405 0.43 ;
      RECT 477.635 0.17 477.895 11.5 ;
      RECT 478.145 0.17 478.405 11.5 ;
      RECT 477.16 118.025 477.36 118.755 ;
      RECT 477.655 118.025 477.855 118.755 ;
      RECT 478.655 0.17 479.425 0.94 ;
      RECT 478.655 0.17 478.915 12.9 ;
      RECT 479.165 0.17 479.425 12.9 ;
      RECT 478.155 118.025 478.355 118.755 ;
      RECT 478.655 118.025 478.855 118.755 ;
      RECT 479.15 118.025 479.35 118.755 ;
      RECT 479.675 0.52 479.935 5.815 ;
      RECT 480.53 0.52 480.79 5.16 ;
      RECT 480.53 4.9 481.31 5.16 ;
      RECT 481.05 4.9 481.31 6.64 ;
      RECT 479.97 118.025 480.17 118.755 ;
      RECT 480.465 118.025 480.665 118.755 ;
      RECT 480.965 118.025 481.165 118.755 ;
      RECT 481.465 118.025 481.665 118.755 ;
      RECT 481.96 118.025 482.16 118.755 ;
      RECT 482.78 118.025 482.98 118.755 ;
      RECT 483.275 118.025 483.475 118.755 ;
      RECT 483.775 118.025 483.975 118.755 ;
      RECT 483.93 0.52 484.19 2.335 ;
      RECT 484.275 118.025 484.475 118.755 ;
      RECT 484.44 0.52 484.7 14.11 ;
      RECT 484.77 118.025 484.97 118.755 ;
      RECT 485.815 0.17 486.585 0.94 ;
      RECT 486.325 0.17 486.585 8.7 ;
      RECT 485.815 0.17 486.075 12.9 ;
      RECT 485.305 0.52 485.565 2.485 ;
      RECT 485.59 118.025 485.79 118.755 ;
      RECT 486.835 0.17 487.605 0.43 ;
      RECT 487.345 0.17 487.605 10.48 ;
      RECT 486.835 0.17 487.095 10.99 ;
      RECT 486.085 118.025 486.285 118.755 ;
      RECT 486.585 118.025 486.785 118.755 ;
      RECT 487.085 118.025 487.285 118.755 ;
      RECT 487.58 118.025 487.78 118.755 ;
      RECT 488.875 0.17 489.645 0.43 ;
      RECT 488.875 0.17 489.135 11.5 ;
      RECT 489.385 0.17 489.645 11.5 ;
      RECT 488.4 118.025 488.6 118.755 ;
      RECT 488.895 118.025 489.095 118.755 ;
      RECT 489.895 0.17 490.665 0.94 ;
      RECT 489.895 0.17 490.155 12.9 ;
      RECT 490.405 0.17 490.665 12.9 ;
      RECT 489.395 118.025 489.595 118.755 ;
      RECT 489.895 118.025 490.095 118.755 ;
      RECT 490.39 118.025 490.59 118.755 ;
      RECT 490.915 0.52 491.175 5.815 ;
      RECT 491.77 0.52 492.03 5.16 ;
      RECT 491.77 4.9 492.55 5.16 ;
      RECT 492.29 4.9 492.55 6.64 ;
      RECT 491.21 118.025 491.41 118.755 ;
      RECT 491.705 118.025 491.905 118.755 ;
      RECT 492.205 118.025 492.405 118.755 ;
      RECT 492.705 118.025 492.905 118.755 ;
      RECT 493.2 118.025 493.4 118.755 ;
      RECT 494.02 118.025 494.22 118.755 ;
      RECT 494.515 118.025 494.715 118.755 ;
      RECT 495.015 118.025 495.215 118.755 ;
      RECT 495.17 0.52 495.43 2.335 ;
      RECT 495.515 118.025 495.715 118.755 ;
      RECT 495.68 0.52 495.94 14.11 ;
      RECT 496.01 118.025 496.21 118.755 ;
      RECT 497.055 0.17 497.825 0.94 ;
      RECT 497.565 0.17 497.825 8.7 ;
      RECT 497.055 0.17 497.315 12.9 ;
      RECT 496.545 0.52 496.805 2.485 ;
      RECT 496.83 118.025 497.03 118.755 ;
      RECT 498.075 0.17 498.845 0.43 ;
      RECT 498.585 0.17 498.845 10.48 ;
      RECT 498.075 0.17 498.335 10.99 ;
      RECT 497.325 118.025 497.525 118.755 ;
      RECT 497.825 118.025 498.025 118.755 ;
      RECT 498.325 118.025 498.525 118.755 ;
      RECT 498.82 118.025 499.02 118.755 ;
      RECT 500.115 0.17 500.885 0.43 ;
      RECT 500.115 0.17 500.375 11.5 ;
      RECT 500.625 0.17 500.885 11.5 ;
      RECT 499.64 118.025 499.84 118.755 ;
      RECT 500.135 118.025 500.335 118.755 ;
      RECT 501.135 0.17 501.905 0.94 ;
      RECT 501.135 0.17 501.395 12.9 ;
      RECT 501.645 0.17 501.905 12.9 ;
      RECT 500.635 118.025 500.835 118.755 ;
      RECT 501.135 118.025 501.335 118.755 ;
      RECT 501.63 118.025 501.83 118.755 ;
      RECT 502.155 0.52 502.415 5.815 ;
      RECT 503.01 0.52 503.27 5.16 ;
      RECT 503.01 4.9 503.79 5.16 ;
      RECT 503.53 4.9 503.79 6.64 ;
      RECT 502.45 118.025 502.65 118.755 ;
      RECT 502.945 118.025 503.145 118.755 ;
      RECT 503.445 118.025 503.645 118.755 ;
      RECT 503.945 118.025 504.145 118.755 ;
      RECT 504.44 118.025 504.64 118.755 ;
      RECT 505.26 118.025 505.46 118.755 ;
      RECT 505.755 118.025 505.955 118.755 ;
      RECT 506.255 118.025 506.455 118.755 ;
      RECT 506.41 0.52 506.67 2.335 ;
      RECT 506.755 118.025 506.955 118.755 ;
      RECT 506.92 0.52 507.18 14.11 ;
      RECT 507.25 118.025 507.45 118.755 ;
      RECT 508.295 0.17 509.065 0.94 ;
      RECT 508.805 0.17 509.065 8.7 ;
      RECT 508.295 0.17 508.555 12.9 ;
      RECT 507.785 0.52 508.045 2.485 ;
      RECT 508.07 118.025 508.27 118.755 ;
      RECT 509.315 0.17 510.085 0.43 ;
      RECT 509.825 0.17 510.085 10.48 ;
      RECT 509.315 0.17 509.575 10.99 ;
      RECT 508.565 118.025 508.765 118.755 ;
      RECT 509.065 118.025 509.265 118.755 ;
      RECT 509.565 118.025 509.765 118.755 ;
      RECT 510.06 118.025 510.26 118.755 ;
      RECT 511.355 0.17 512.125 0.43 ;
      RECT 511.355 0.17 511.615 11.5 ;
      RECT 511.865 0.17 512.125 11.5 ;
      RECT 510.88 118.025 511.08 118.755 ;
      RECT 511.375 118.025 511.575 118.755 ;
      RECT 512.375 0.17 513.145 0.94 ;
      RECT 512.375 0.17 512.635 12.9 ;
      RECT 512.885 0.17 513.145 12.9 ;
      RECT 511.875 118.025 512.075 118.755 ;
      RECT 512.375 118.025 512.575 118.755 ;
      RECT 512.87 118.025 513.07 118.755 ;
      RECT 513.395 0.52 513.655 5.815 ;
      RECT 514.25 0.52 514.51 5.16 ;
      RECT 514.25 4.9 515.03 5.16 ;
      RECT 514.77 4.9 515.03 6.64 ;
      RECT 513.69 118.025 513.89 118.755 ;
      RECT 514.185 118.025 514.385 118.755 ;
      RECT 514.685 118.025 514.885 118.755 ;
      RECT 515.185 118.025 515.385 118.755 ;
      RECT 515.68 118.025 515.88 118.755 ;
      RECT 516.5 118.025 516.7 118.755 ;
      RECT 516.995 118.025 517.195 118.755 ;
      RECT 517.495 118.025 517.695 118.755 ;
      RECT 517.65 0.52 517.91 2.335 ;
      RECT 517.995 118.025 518.195 118.755 ;
      RECT 518.16 0.52 518.42 14.11 ;
      RECT 518.49 118.025 518.69 118.755 ;
      RECT 519.535 0.17 520.305 0.94 ;
      RECT 520.045 0.17 520.305 8.7 ;
      RECT 519.535 0.17 519.795 12.9 ;
      RECT 519.025 0.52 519.285 2.485 ;
      RECT 519.31 118.025 519.51 118.755 ;
      RECT 520.555 0.17 521.325 0.43 ;
      RECT 521.065 0.17 521.325 10.48 ;
      RECT 520.555 0.17 520.815 10.99 ;
      RECT 519.805 118.025 520.005 118.755 ;
      RECT 520.305 118.025 520.505 118.755 ;
      RECT 520.805 118.025 521.005 118.755 ;
      RECT 521.3 118.025 521.5 118.755 ;
      RECT 522.595 0.17 523.365 0.43 ;
      RECT 522.595 0.17 522.855 11.5 ;
      RECT 523.105 0.17 523.365 11.5 ;
      RECT 522.12 118.025 522.32 118.755 ;
      RECT 522.615 118.025 522.815 118.755 ;
      RECT 523.615 0.17 524.385 0.94 ;
      RECT 523.615 0.17 523.875 12.9 ;
      RECT 524.125 0.17 524.385 12.9 ;
      RECT 523.115 118.025 523.315 118.755 ;
      RECT 523.615 118.025 523.815 118.755 ;
      RECT 524.11 118.025 524.31 118.755 ;
      RECT 524.635 0.52 524.895 5.815 ;
      RECT 525.49 0.52 525.75 5.16 ;
      RECT 525.49 4.9 526.27 5.16 ;
      RECT 526.01 4.9 526.27 6.64 ;
      RECT 524.93 118.025 525.13 118.755 ;
      RECT 525.425 118.025 525.625 118.755 ;
      RECT 525.925 118.025 526.125 118.755 ;
      RECT 526.425 118.025 526.625 118.755 ;
      RECT 526.92 118.025 527.12 118.755 ;
      RECT 527.74 118.025 527.94 118.755 ;
      RECT 528.235 118.025 528.435 118.755 ;
      RECT 528.735 118.025 528.935 118.755 ;
      RECT 528.89 0.52 529.15 2.335 ;
      RECT 529.235 118.025 529.435 118.755 ;
      RECT 529.4 0.52 529.66 14.11 ;
      RECT 529.73 118.025 529.93 118.755 ;
      RECT 530.775 0.17 531.545 0.94 ;
      RECT 531.285 0.17 531.545 8.7 ;
      RECT 530.775 0.17 531.035 12.9 ;
      RECT 530.265 0.52 530.525 2.485 ;
      RECT 530.55 118.025 530.75 118.755 ;
      RECT 531.795 0.17 532.565 0.43 ;
      RECT 532.305 0.17 532.565 10.48 ;
      RECT 531.795 0.17 532.055 10.99 ;
      RECT 531.045 118.025 531.245 118.755 ;
      RECT 531.545 118.025 531.745 118.755 ;
      RECT 532.045 118.025 532.245 118.755 ;
      RECT 532.54 118.025 532.74 118.755 ;
      RECT 533.835 0.17 534.605 0.43 ;
      RECT 533.835 0.17 534.095 11.5 ;
      RECT 534.345 0.17 534.605 11.5 ;
      RECT 533.36 118.025 533.56 118.755 ;
      RECT 533.855 118.025 534.055 118.755 ;
      RECT 534.855 0.17 535.625 0.94 ;
      RECT 534.855 0.17 535.115 12.9 ;
      RECT 535.365 0.17 535.625 12.9 ;
      RECT 534.355 118.025 534.555 118.755 ;
      RECT 534.855 118.025 535.055 118.755 ;
      RECT 535.35 118.025 535.55 118.755 ;
      RECT 535.875 0.52 536.135 5.815 ;
      RECT 536.73 0.52 536.99 5.16 ;
      RECT 536.73 4.9 537.51 5.16 ;
      RECT 537.25 4.9 537.51 6.64 ;
      RECT 536.17 118.025 536.37 118.755 ;
      RECT 536.665 118.025 536.865 118.755 ;
      RECT 537.165 118.025 537.365 118.755 ;
      RECT 537.665 118.025 537.865 118.755 ;
      RECT 538.16 118.025 538.36 118.755 ;
      RECT 538.98 118.025 539.18 118.755 ;
      RECT 539.475 118.025 539.675 118.755 ;
      RECT 539.975 118.025 540.175 118.755 ;
      RECT 540.13 0.52 540.39 2.335 ;
      RECT 540.475 118.025 540.675 118.755 ;
      RECT 540.64 0.52 540.9 14.11 ;
      RECT 540.97 118.025 541.17 118.755 ;
      RECT 542.015 0.17 542.785 0.94 ;
      RECT 542.525 0.17 542.785 8.7 ;
      RECT 542.015 0.17 542.275 12.9 ;
      RECT 541.505 0.52 541.765 2.485 ;
      RECT 541.79 118.025 541.99 118.755 ;
      RECT 543.035 0.17 543.805 0.43 ;
      RECT 543.545 0.17 543.805 10.48 ;
      RECT 543.035 0.17 543.295 10.99 ;
      RECT 542.285 118.025 542.485 118.755 ;
      RECT 542.785 118.025 542.985 118.755 ;
      RECT 543.285 118.025 543.485 118.755 ;
      RECT 543.78 118.025 543.98 118.755 ;
      RECT 545.075 0.17 545.845 0.43 ;
      RECT 545.075 0.17 545.335 11.5 ;
      RECT 545.585 0.17 545.845 11.5 ;
      RECT 544.6 118.025 544.8 118.755 ;
      RECT 545.095 118.025 545.295 118.755 ;
      RECT 546.095 0.17 546.865 0.94 ;
      RECT 546.095 0.17 546.355 12.9 ;
      RECT 546.605 0.17 546.865 12.9 ;
      RECT 545.595 118.025 545.795 118.755 ;
      RECT 546.095 118.025 546.295 118.755 ;
      RECT 546.59 118.025 546.79 118.755 ;
      RECT 547.115 0.52 547.375 5.815 ;
      RECT 547.97 0.52 548.23 5.16 ;
      RECT 547.97 4.9 548.75 5.16 ;
      RECT 548.49 4.9 548.75 6.64 ;
      RECT 547.41 118.025 547.61 118.755 ;
      RECT 547.905 118.025 548.105 118.755 ;
      RECT 548.405 118.025 548.605 118.755 ;
      RECT 548.905 118.025 549.105 118.755 ;
      RECT 549.4 118.025 549.6 118.755 ;
      RECT 550.22 118.025 550.42 118.755 ;
      RECT 550.715 118.025 550.915 118.755 ;
      RECT 551.215 118.025 551.415 118.755 ;
      RECT 551.37 0.52 551.63 2.335 ;
      RECT 551.715 118.025 551.915 118.755 ;
      RECT 551.88 0.52 552.14 14.11 ;
      RECT 552.21 118.025 552.41 118.755 ;
      RECT 553.255 0.17 554.025 0.94 ;
      RECT 553.765 0.17 554.025 8.7 ;
      RECT 553.255 0.17 553.515 12.9 ;
      RECT 552.745 0.52 553.005 2.485 ;
      RECT 553.03 118.025 553.23 118.755 ;
      RECT 554.275 0.17 555.045 0.43 ;
      RECT 554.785 0.17 555.045 10.48 ;
      RECT 554.275 0.17 554.535 10.99 ;
      RECT 553.525 118.025 553.725 118.755 ;
      RECT 554.025 118.025 554.225 118.755 ;
      RECT 554.525 118.025 554.725 118.755 ;
      RECT 555.02 118.025 555.22 118.755 ;
      RECT 556.315 0.17 557.085 0.43 ;
      RECT 556.315 0.17 556.575 11.5 ;
      RECT 556.825 0.17 557.085 11.5 ;
      RECT 555.84 118.025 556.04 118.755 ;
      RECT 556.335 118.025 556.535 118.755 ;
      RECT 557.335 0.17 558.105 0.94 ;
      RECT 557.335 0.17 557.595 12.9 ;
      RECT 557.845 0.17 558.105 12.9 ;
      RECT 556.835 118.025 557.035 118.755 ;
      RECT 557.335 118.025 557.535 118.755 ;
      RECT 557.83 118.025 558.03 118.755 ;
      RECT 558.355 0.52 558.615 5.815 ;
      RECT 559.21 0.52 559.47 5.16 ;
      RECT 559.21 4.9 559.99 5.16 ;
      RECT 559.73 4.9 559.99 6.64 ;
      RECT 558.65 118.025 558.85 118.755 ;
      RECT 559.145 118.025 559.345 118.755 ;
      RECT 559.645 118.025 559.845 118.755 ;
      RECT 560.145 118.025 560.345 118.755 ;
      RECT 560.64 118.025 560.84 118.755 ;
      RECT 561.46 118.025 561.66 118.755 ;
      RECT 561.955 118.025 562.155 118.755 ;
      RECT 562.455 118.025 562.655 118.755 ;
      RECT 562.61 0.52 562.87 2.335 ;
      RECT 562.955 118.025 563.155 118.755 ;
      RECT 563.12 0.52 563.38 14.11 ;
      RECT 563.45 118.025 563.65 118.755 ;
      RECT 564.495 0.17 565.265 0.94 ;
      RECT 565.005 0.17 565.265 8.7 ;
      RECT 564.495 0.17 564.755 12.9 ;
      RECT 563.985 0.52 564.245 2.485 ;
      RECT 564.27 118.025 564.47 118.755 ;
      RECT 565.515 0.17 566.285 0.43 ;
      RECT 566.025 0.17 566.285 10.48 ;
      RECT 565.515 0.17 565.775 10.99 ;
      RECT 564.765 118.025 564.965 118.755 ;
      RECT 565.265 118.025 565.465 118.755 ;
      RECT 565.765 118.025 565.965 118.755 ;
      RECT 566.26 118.025 566.46 118.755 ;
      RECT 567.555 0.17 568.325 0.43 ;
      RECT 567.555 0.17 567.815 11.5 ;
      RECT 568.065 0.17 568.325 11.5 ;
      RECT 567.08 118.025 567.28 118.755 ;
      RECT 567.575 118.025 567.775 118.755 ;
      RECT 568.575 0.17 569.345 0.94 ;
      RECT 568.575 0.17 568.835 12.9 ;
      RECT 569.085 0.17 569.345 12.9 ;
      RECT 568.075 118.025 568.275 118.755 ;
      RECT 568.575 118.025 568.775 118.755 ;
      RECT 569.07 118.025 569.27 118.755 ;
      RECT 569.595 0.52 569.855 5.815 ;
      RECT 570.45 0.52 570.71 5.16 ;
      RECT 570.45 4.9 571.23 5.16 ;
      RECT 570.97 4.9 571.23 6.64 ;
      RECT 569.89 118.025 570.09 118.755 ;
      RECT 570.385 118.025 570.585 118.755 ;
      RECT 570.885 118.025 571.085 118.755 ;
      RECT 571.385 118.025 571.585 118.755 ;
      RECT 571.88 118.025 572.08 118.755 ;
      RECT 572.7 118.025 572.9 118.755 ;
      RECT 573.195 118.025 573.395 118.755 ;
      RECT 573.695 118.025 573.895 118.755 ;
      RECT 573.85 0.52 574.11 2.335 ;
      RECT 574.195 118.025 574.395 118.755 ;
      RECT 574.36 0.52 574.62 14.11 ;
      RECT 574.69 118.025 574.89 118.755 ;
      RECT 575.735 0.17 576.505 0.94 ;
      RECT 576.245 0.17 576.505 8.7 ;
      RECT 575.735 0.17 575.995 12.9 ;
      RECT 575.225 0.52 575.485 2.485 ;
      RECT 575.51 118.025 575.71 118.755 ;
      RECT 576.755 0.17 577.525 0.43 ;
      RECT 577.265 0.17 577.525 10.48 ;
      RECT 576.755 0.17 577.015 10.99 ;
      RECT 576.005 118.025 576.205 118.755 ;
      RECT 576.505 118.025 576.705 118.755 ;
      RECT 577.005 118.025 577.205 118.755 ;
      RECT 577.5 118.025 577.7 118.755 ;
      RECT 578.795 0.17 579.565 0.43 ;
      RECT 578.795 0.17 579.055 11.5 ;
      RECT 579.305 0.17 579.565 11.5 ;
      RECT 578.32 118.025 578.52 118.755 ;
      RECT 578.815 118.025 579.015 118.755 ;
      RECT 579.815 0.17 580.585 0.94 ;
      RECT 579.815 0.17 580.075 12.9 ;
      RECT 580.325 0.17 580.585 12.9 ;
      RECT 579.315 118.025 579.515 118.755 ;
      RECT 579.815 118.025 580.015 118.755 ;
      RECT 580.31 118.025 580.51 118.755 ;
      RECT 580.835 0.52 581.095 5.815 ;
      RECT 581.69 0.52 581.95 5.16 ;
      RECT 581.69 4.9 582.47 5.16 ;
      RECT 582.21 4.9 582.47 6.64 ;
      RECT 581.13 118.025 581.33 118.755 ;
      RECT 581.625 118.025 581.825 118.755 ;
      RECT 582.125 118.025 582.325 118.755 ;
      RECT 582.625 118.025 582.825 118.755 ;
      RECT 583.12 118.025 583.32 118.755 ;
      RECT 583.94 118.025 584.14 118.755 ;
      RECT 584.435 118.025 584.635 118.755 ;
      RECT 584.935 118.025 585.135 118.755 ;
      RECT 585.09 0.52 585.35 2.335 ;
      RECT 585.435 118.025 585.635 118.755 ;
      RECT 585.6 0.52 585.86 14.11 ;
      RECT 585.93 118.025 586.13 118.755 ;
      RECT 586.975 0.17 587.745 0.94 ;
      RECT 587.485 0.17 587.745 8.7 ;
      RECT 586.975 0.17 587.235 12.9 ;
      RECT 586.465 0.52 586.725 2.485 ;
      RECT 586.75 118.025 586.95 118.755 ;
      RECT 587.995 0.17 588.765 0.43 ;
      RECT 588.505 0.17 588.765 10.48 ;
      RECT 587.995 0.17 588.255 10.99 ;
      RECT 587.245 118.025 587.445 118.755 ;
      RECT 587.745 118.025 587.945 118.755 ;
      RECT 588.245 118.025 588.445 118.755 ;
      RECT 588.74 118.025 588.94 118.755 ;
      RECT 590.035 0.17 590.805 0.43 ;
      RECT 590.035 0.17 590.295 11.5 ;
      RECT 590.545 0.17 590.805 11.5 ;
      RECT 589.56 118.025 589.76 118.755 ;
      RECT 590.055 118.025 590.255 118.755 ;
      RECT 591.055 0.17 591.825 0.94 ;
      RECT 591.055 0.17 591.315 12.9 ;
      RECT 591.565 0.17 591.825 12.9 ;
      RECT 590.555 118.025 590.755 118.755 ;
      RECT 591.055 118.025 591.255 118.755 ;
      RECT 591.55 118.025 591.75 118.755 ;
      RECT 592.075 0.52 592.335 5.815 ;
      RECT 592.93 0.52 593.19 5.16 ;
      RECT 592.93 4.9 593.71 5.16 ;
      RECT 593.45 4.9 593.71 6.64 ;
      RECT 592.37 118.025 592.57 118.755 ;
      RECT 592.865 118.025 593.065 118.755 ;
      RECT 593.365 118.025 593.565 118.755 ;
      RECT 593.865 118.025 594.065 118.755 ;
      RECT 594.36 118.025 594.56 118.755 ;
      RECT 595.18 118.025 595.38 118.755 ;
      RECT 596.175 45.465 596.375 118.755 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 184.505 0 189.335 118.78 ;
      RECT 195.745 0 200.575 118.78 ;
      RECT 206.985 0 211.815 118.78 ;
      RECT 218.225 0 223.055 118.78 ;
      RECT 229.465 0 234.295 118.78 ;
      RECT 240.705 0 245.535 118.78 ;
      RECT 251.945 0 256.775 118.78 ;
      RECT 263.185 0 268.015 118.78 ;
      RECT 284.24 0 290.61 118.78 ;
      RECT 299.55 0 300.81 118.78 ;
      RECT 328.465 0 333.295 118.78 ;
      RECT 339.705 0 344.535 118.78 ;
      RECT 350.945 0 355.775 118.78 ;
      RECT 362.185 0 367.015 118.78 ;
      RECT 373.425 0 378.255 118.78 ;
      RECT 384.665 0 389.495 118.78 ;
      RECT 395.905 0 400.735 118.78 ;
      RECT 407.145 0 411.975 118.78 ;
      RECT 418.385 0 423.215 118.78 ;
      RECT 429.625 0 434.455 118.78 ;
      RECT 440.865 0 445.695 118.78 ;
      RECT 452.105 0 456.935 118.78 ;
      RECT 463.345 0 468.175 118.78 ;
      RECT 474.585 0 479.415 118.78 ;
      RECT 485.825 0 490.655 118.78 ;
      RECT 497.065 0 501.895 118.78 ;
      RECT 508.305 0 513.135 118.78 ;
      RECT 519.545 0 524.375 118.78 ;
      RECT 530.785 0 535.615 118.78 ;
      RECT 542.025 0 546.855 118.78 ;
      RECT 553.265 0 558.095 118.78 ;
      RECT 564.505 0 569.335 118.78 ;
      RECT 575.745 0 580.575 118.78 ;
      RECT 586.985 0 591.815 118.78 ;
      RECT 291.9 0 292.14 118.78 ;
      RECT 293.43 0 293.67 118.78 ;
      RECT 296.49 0 296.73 118.78 ;
      RECT 298.02 0 298.26 118.78 ;
      RECT 305.15 0 314.07 118.78 ;
      RECT 0 0 3.03 118.78 ;
      RECT 4.655 0.17 9.505 118.78 ;
      RECT 11.65 0 14.27 118.78 ;
      RECT 15.895 0.17 20.745 118.78 ;
      RECT 22.89 0 25.51 118.78 ;
      RECT 27.135 0.17 31.985 118.78 ;
      RECT 34.13 0 36.75 118.78 ;
      RECT 38.375 0.17 43.225 118.78 ;
      RECT 45.37 0 47.99 118.78 ;
      RECT 49.615 0.17 54.465 118.78 ;
      RECT 56.61 0 59.23 118.78 ;
      RECT 60.855 0.17 65.705 118.78 ;
      RECT 67.85 0 70.47 118.78 ;
      RECT 72.095 0.17 76.945 118.78 ;
      RECT 79.09 0 81.71 118.78 ;
      RECT 83.335 0.17 88.185 118.78 ;
      RECT 90.33 0 92.95 118.78 ;
      RECT 94.575 0.17 99.425 118.78 ;
      RECT 101.57 0 104.19 118.78 ;
      RECT 105.815 0.17 110.665 118.78 ;
      RECT 112.81 0 115.43 118.78 ;
      RECT 117.055 0.17 121.905 118.78 ;
      RECT 124.05 0 126.67 118.78 ;
      RECT 128.295 0.17 133.145 118.78 ;
      RECT 135.29 0 137.91 118.78 ;
      RECT 139.535 0.17 144.385 118.78 ;
      RECT 146.53 0 149.15 118.78 ;
      RECT 150.775 0.17 155.625 118.78 ;
      RECT 157.77 0 160.39 118.78 ;
      RECT 162.015 0.17 166.865 118.78 ;
      RECT 169.01 0 171.63 118.78 ;
      RECT 173.255 0.17 178.105 118.78 ;
      RECT 180.25 0 182.87 118.78 ;
      RECT 184.495 0.17 189.345 118.78 ;
      RECT 191.49 0 194.11 118.78 ;
      RECT 195.735 0.17 200.585 118.78 ;
      RECT 202.73 0 205.35 118.78 ;
      RECT 206.975 0.17 211.825 118.78 ;
      RECT 213.97 0 216.59 118.78 ;
      RECT 218.215 0.17 223.065 118.78 ;
      RECT 225.21 0 227.83 118.78 ;
      RECT 229.455 0.17 234.305 118.78 ;
      RECT 236.45 0 239.07 118.78 ;
      RECT 240.695 0.17 245.545 118.78 ;
      RECT 247.69 0 250.31 118.78 ;
      RECT 251.935 0.17 256.785 118.78 ;
      RECT 258.93 0 261.55 118.78 ;
      RECT 263.175 0.17 268.025 118.78 ;
      RECT 270.17 0 281.95 118.78 ;
      RECT 284.24 0.17 290.62 118.78 ;
      RECT 291.89 0.3 292.15 118.78 ;
      RECT 293.42 0.3 293.68 118.78 ;
      RECT 296.48 0.3 296.74 118.78 ;
      RECT 298.01 0.3 298.27 118.78 ;
      RECT 299.55 0.17 300.82 118.78 ;
      RECT 299.54 0.3 300.82 118.78 ;
      RECT 305.15 0.3 314.08 118.78 ;
      RECT 314.85 0 326.31 118.78 ;
      RECT 314.84 0.17 326.31 118.78 ;
      RECT 328.455 0.17 333.305 118.78 ;
      RECT 334.93 0 337.55 118.78 ;
      RECT 339.695 0.17 344.545 118.78 ;
      RECT 346.17 0 348.79 118.78 ;
      RECT 350.935 0.17 355.785 118.78 ;
      RECT 357.41 0 360.03 118.78 ;
      RECT 362.175 0.17 367.025 118.78 ;
      RECT 368.65 0 371.27 118.78 ;
      RECT 373.415 0.17 378.265 118.78 ;
      RECT 379.89 0 382.51 118.78 ;
      RECT 384.655 0.17 389.505 118.78 ;
      RECT 391.13 0 393.75 118.78 ;
      RECT 395.895 0.17 400.745 118.78 ;
      RECT 402.37 0 404.99 118.78 ;
      RECT 407.135 0.17 411.985 118.78 ;
      RECT 413.61 0 416.23 118.78 ;
      RECT 418.375 0.17 423.225 118.78 ;
      RECT 424.85 0 427.47 118.78 ;
      RECT 429.615 0.17 434.465 118.78 ;
      RECT 436.09 0 438.71 118.78 ;
      RECT 440.855 0.17 445.705 118.78 ;
      RECT 447.33 0 449.95 118.78 ;
      RECT 452.095 0.17 456.945 118.78 ;
      RECT 458.57 0 461.19 118.78 ;
      RECT 463.335 0.17 468.185 118.78 ;
      RECT 469.81 0 472.43 118.78 ;
      RECT 474.575 0.17 479.425 118.78 ;
      RECT 481.05 0 483.67 118.78 ;
      RECT 485.815 0.17 490.665 118.78 ;
      RECT 492.29 0 494.91 118.78 ;
      RECT 497.055 0.17 501.905 118.78 ;
      RECT 503.53 0 506.15 118.78 ;
      RECT 508.295 0.17 513.145 118.78 ;
      RECT 514.77 0 517.39 118.78 ;
      RECT 519.535 0.17 524.385 118.78 ;
      RECT 526.01 0 528.63 118.78 ;
      RECT 530.775 0.17 535.625 118.78 ;
      RECT 537.25 0 539.87 118.78 ;
      RECT 542.015 0.17 546.865 118.78 ;
      RECT 548.49 0 551.11 118.78 ;
      RECT 553.255 0.17 558.105 118.78 ;
      RECT 559.73 0 562.35 118.78 ;
      RECT 564.495 0.17 569.345 118.78 ;
      RECT 570.97 0 573.59 118.78 ;
      RECT 575.735 0.17 580.585 118.78 ;
      RECT 582.21 0 584.83 118.78 ;
      RECT 586.975 0.17 591.825 118.78 ;
      RECT 593.45 0 596.48 118.78 ;
      RECT 0 0.52 596.48 118.78 ;
      RECT 4.665 0 9.495 118.78 ;
      RECT 15.905 0 20.735 118.78 ;
      RECT 27.145 0 31.975 118.78 ;
      RECT 38.385 0 43.215 118.78 ;
      RECT 49.625 0 54.455 118.78 ;
      RECT 60.865 0 65.695 118.78 ;
      RECT 72.105 0 76.935 118.78 ;
      RECT 83.345 0 88.175 118.78 ;
      RECT 94.585 0 99.415 118.78 ;
      RECT 105.825 0 110.655 118.78 ;
      RECT 117.065 0 121.895 118.78 ;
      RECT 128.305 0 133.135 118.78 ;
      RECT 139.545 0 144.375 118.78 ;
      RECT 150.785 0 155.615 118.78 ;
      RECT 162.025 0 166.855 118.78 ;
      RECT 173.265 0 178.095 118.78 ;
    LAYER Metal3 ;
      RECT 0 0 596.48 118.78 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 0 39.085 9.62 45.205 ;
      RECT 0 0 4 118.78 ;
      RECT 7.33 0 9.62 118.78 ;
      RECT 12.95 39.085 20.86 45.205 ;
      RECT 12.95 0 15.24 118.78 ;
      RECT 18.57 0 20.86 118.78 ;
      RECT 24.19 39.085 32.1 45.205 ;
      RECT 24.19 0 26.48 118.78 ;
      RECT 29.81 0 32.1 118.78 ;
      RECT 35.43 39.085 43.34 45.205 ;
      RECT 35.43 0 37.72 118.78 ;
      RECT 41.05 0 43.34 118.78 ;
      RECT 46.67 39.085 54.58 45.205 ;
      RECT 46.67 0 48.96 118.78 ;
      RECT 52.29 0 54.58 118.78 ;
      RECT 57.91 39.085 65.82 45.205 ;
      RECT 57.91 0 60.2 118.78 ;
      RECT 63.53 0 65.82 118.78 ;
      RECT 69.15 39.085 77.06 45.205 ;
      RECT 69.15 0 71.44 118.78 ;
      RECT 74.77 0 77.06 118.78 ;
      RECT 80.39 39.085 88.3 45.205 ;
      RECT 80.39 0 82.68 118.78 ;
      RECT 86.01 0 88.3 118.78 ;
      RECT 91.63 39.085 99.54 45.205 ;
      RECT 91.63 0 93.92 118.78 ;
      RECT 97.25 0 99.54 118.78 ;
      RECT 102.87 39.085 110.78 45.205 ;
      RECT 102.87 0 105.16 118.78 ;
      RECT 108.49 0 110.78 118.78 ;
      RECT 114.11 39.085 122.02 45.205 ;
      RECT 114.11 0 116.4 118.78 ;
      RECT 119.73 0 122.02 118.78 ;
      RECT 125.35 39.085 133.26 45.205 ;
      RECT 125.35 0 127.64 118.78 ;
      RECT 130.97 0 133.26 118.78 ;
      RECT 136.59 39.085 144.5 45.205 ;
      RECT 136.59 0 138.88 118.78 ;
      RECT 142.21 0 144.5 118.78 ;
      RECT 147.83 39.085 155.74 45.205 ;
      RECT 147.83 0 150.12 118.78 ;
      RECT 153.45 0 155.74 118.78 ;
      RECT 159.07 39.085 166.98 45.205 ;
      RECT 159.07 0 161.36 118.78 ;
      RECT 164.69 0 166.98 118.78 ;
      RECT 170.31 39.085 178.22 45.205 ;
      RECT 170.31 0 172.6 118.78 ;
      RECT 175.93 0 178.22 118.78 ;
      RECT 181.55 39.085 189.46 45.205 ;
      RECT 181.55 0 183.84 118.78 ;
      RECT 187.17 0 189.46 118.78 ;
      RECT 192.79 39.085 200.7 45.205 ;
      RECT 192.79 0 195.08 118.78 ;
      RECT 198.41 0 200.7 118.78 ;
      RECT 204.03 39.085 211.94 45.205 ;
      RECT 204.03 0 206.32 118.78 ;
      RECT 209.65 0 211.94 118.78 ;
      RECT 215.27 39.085 223.18 45.205 ;
      RECT 215.27 0 217.56 118.78 ;
      RECT 220.89 0 223.18 118.78 ;
      RECT 226.51 39.085 234.42 45.205 ;
      RECT 226.51 0 228.8 118.78 ;
      RECT 232.13 0 234.42 118.78 ;
      RECT 237.75 39.085 245.66 45.205 ;
      RECT 237.75 0 240.04 118.78 ;
      RECT 243.37 0 245.66 118.78 ;
      RECT 248.99 39.085 256.9 45.205 ;
      RECT 248.99 0 251.28 118.78 ;
      RECT 254.61 0 256.9 118.78 ;
      RECT 260.23 39.085 268.14 45.205 ;
      RECT 260.23 0 262.52 118.78 ;
      RECT 265.85 0 268.14 118.78 ;
      RECT 271.47 0 278.55 118.78 ;
      RECT 281.88 0 283.7 118.78 ;
      RECT 287.03 0 288.85 118.78 ;
      RECT 292.18 0 294 118.78 ;
      RECT 297.33 0 299.15 118.78 ;
      RECT 302.48 0 304.3 118.78 ;
      RECT 328.34 39.085 336.25 45.205 ;
      RECT 328.34 0 330.63 118.78 ;
      RECT 333.96 0 336.25 118.78 ;
      RECT 339.58 39.085 347.49 45.205 ;
      RECT 339.58 0 341.87 118.78 ;
      RECT 345.2 0 347.49 118.78 ;
      RECT 350.82 39.085 358.73 45.205 ;
      RECT 350.82 0 353.11 118.78 ;
      RECT 356.44 0 358.73 118.78 ;
      RECT 362.06 39.085 369.97 45.205 ;
      RECT 362.06 0 364.35 118.78 ;
      RECT 367.68 0 369.97 118.78 ;
      RECT 373.3 39.085 381.21 45.205 ;
      RECT 373.3 0 375.59 118.78 ;
      RECT 378.92 0 381.21 118.78 ;
      RECT 384.54 39.085 392.45 45.205 ;
      RECT 384.54 0 386.83 118.78 ;
      RECT 390.16 0 392.45 118.78 ;
      RECT 395.78 39.085 403.69 45.205 ;
      RECT 395.78 0 398.07 118.78 ;
      RECT 401.4 0 403.69 118.78 ;
      RECT 407.02 39.085 414.93 45.205 ;
      RECT 407.02 0 409.31 118.78 ;
      RECT 412.64 0 414.93 118.78 ;
      RECT 418.26 39.085 426.17 45.205 ;
      RECT 418.26 0 420.55 118.78 ;
      RECT 423.88 0 426.17 118.78 ;
      RECT 429.5 39.085 437.41 45.205 ;
      RECT 429.5 0 431.79 118.78 ;
      RECT 435.12 0 437.41 118.78 ;
      RECT 440.74 39.085 448.65 45.205 ;
      RECT 440.74 0 443.03 118.78 ;
      RECT 446.36 0 448.65 118.78 ;
      RECT 451.98 39.085 459.89 45.205 ;
      RECT 451.98 0 454.27 118.78 ;
      RECT 457.6 0 459.89 118.78 ;
      RECT 463.22 39.085 471.13 45.205 ;
      RECT 463.22 0 465.51 118.78 ;
      RECT 468.84 0 471.13 118.78 ;
      RECT 474.46 39.085 482.37 45.205 ;
      RECT 474.46 0 476.75 118.78 ;
      RECT 480.08 0 482.37 118.78 ;
      RECT 485.7 39.085 493.61 45.205 ;
      RECT 485.7 0 487.99 118.78 ;
      RECT 491.32 0 493.61 118.78 ;
      RECT 496.94 39.085 504.85 45.205 ;
      RECT 496.94 0 499.23 118.78 ;
      RECT 502.56 0 504.85 118.78 ;
      RECT 508.18 39.085 516.09 45.205 ;
      RECT 508.18 0 510.47 118.78 ;
      RECT 513.8 0 516.09 118.78 ;
      RECT 519.42 39.085 527.33 45.205 ;
      RECT 519.42 0 521.71 118.78 ;
      RECT 525.04 0 527.33 118.78 ;
      RECT 530.66 39.085 538.57 45.205 ;
      RECT 530.66 0 532.95 118.78 ;
      RECT 536.28 0 538.57 118.78 ;
      RECT 541.9 39.085 549.81 45.205 ;
      RECT 541.9 0 544.19 118.78 ;
      RECT 547.52 0 549.81 118.78 ;
      RECT 553.14 39.085 561.05 45.205 ;
      RECT 553.14 0 555.43 118.78 ;
      RECT 558.76 0 561.05 118.78 ;
      RECT 564.38 39.085 572.29 45.205 ;
      RECT 564.38 0 566.67 118.78 ;
      RECT 570 0 572.29 118.78 ;
      RECT 575.62 39.085 583.53 45.205 ;
      RECT 575.62 0 577.91 118.78 ;
      RECT 581.24 0 583.53 118.78 ;
      RECT 586.86 39.085 596.48 45.205 ;
      RECT 586.86 0 589.15 118.78 ;
      RECT 592.48 0 596.48 118.78 ;
      RECT 307.63 0 309.45 118.78 ;
      RECT 312.78 0 314.6 118.78 ;
      RECT 317.93 0 325.01 118.78 ;
  END
END RM_IHPSG13_1P_256x48_c2_bm_bist

END LIBRARY
