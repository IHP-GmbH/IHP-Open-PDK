*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT cap_cmim
C0 PLUS1 MINUS1 cap_cmim w=6.99u l=6.99u m=1
C1 PLUS2 MINUS2 cap_cmim w=6.99u l=6.99u m=2
C2 PLUS3 MINUS3 cap_cmim w=6.99u l=6.99u m=3
.ENDS
