*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT npn13G2v
Q1 net1 net2 net3 sub npn13G2v m=1 le=1.0u  we=120.00n
Q2 net4 net5 net6 sub npn13G2v m=1 le=1.15u we=120.00n
Q3 net7 net8 net9 sub npn13G2v m=2 le=1.0u  we=120.00n

* Extra patterns
Q_pattern_1  c_1  b_1  e_1  sub npn13G2v we=0.12u le=1.63u 
Q_pattern_2  c_2  b_2  e_2  sub npn13G2v we=0.12u le=3.14u 
Q_pattern_3  c_3  b_3  e_3  sub npn13G2v we=0.12u le=4.45u 
Q_pattern_4  c_4  b_4  e_4  sub npn13G2v we=0.12u le=2.17u 
Q_pattern_5  c_5  b_5  e_5  sub npn13G2v we=0.12u le=2.55u 
Q_pattern_6  c_6  b_6  e_6  sub npn13G2v we=0.12u le=3.52u 
Q_pattern_7  c_7  b_7  e_7  sub npn13G2v we=0.12u le=3.22u 
Q_pattern_8  c_8  b_8  e_8  sub npn13G2v we=0.12u le=2.79u 
Q_pattern_9  c_9  b_9  e_9  sub npn13G2v we=0.12u le=2.79u 
Q_pattern_10 c_10 b_10 e_10 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_11 c_11 b_11 e_11 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_12 c_12 b_12 e_12 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_13 c_13 b_13 e_13 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_14 c_14 b_14 e_14 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_15 c_15 b_15 e_15 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_16 c_16 b_16 e_16 sub npn13G2v we=0.12u le=1.63u 
Q_pattern_17 c_17 b_17 e_17 sub npn13G2v we=0.12u le=1.63u 
Q_pattern_18 c_18 b_18 e_18 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_19 c_19 b_19 e_19 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_20 c_20 b_20 e_20 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_21 c_21 b_21 e_21 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_22 c_22 b_22 e_22 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_23 c_23 b_23 e_23 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_24 c_24 b_24 e_24 sub npn13G2v we=0.12u le=2.79u 
Q_pattern_25 c_25 b_25 e_25 sub npn13G2v we=0.12u le=2.79u 
Q_pattern_26 c_26 b_26 e_26 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_27 c_27 b_27 e_27 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_28 c_28 b_28 e_28 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_29 c_29 b_29 e_29 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_30 c_30 b_30 e_30 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_31 c_31 b_31 e_31 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_32 c_32 b_32 e_32 sub npn13G2v we=0.12u le=1.63u 
Q_pattern_33 c_33 b_33 e_33 sub npn13G2v we=0.12u le=1.63u 
Q_pattern_34 c_34 b_34 e_34 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_35 c_35 b_35 e_35 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_36 c_36 b_36 e_36 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_37 c_37 b_37 e_37 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_38 c_38 b_38 e_38 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_39 c_39 b_39 e_39 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_40 c_40 b_40 e_40 sub npn13G2v we=0.12u le=2.79u 
Q_pattern_41 c_41 b_41 e_41 sub npn13G2v we=0.12u le=2.79u 
Q_pattern_42 c_42 b_42 e_42 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_43 c_43 b_43 e_43 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_44 c_44 b_44 e_44 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_45 c_45 b_45 e_45 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_46 c_46 b_46 e_46 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_47 c_47 b_47 e_47 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_48 c_48 b_48 e_48 sub npn13G2v we=0.12u le=1.63u 
Q_pattern_49 c_49 b_49 e_49 sub npn13G2v we=0.12u le=1.63u 
Q_pattern_50 c_50 b_50 e_50 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_51 c_51 b_51 e_51 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_52 c_52 b_52 e_52 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_53 c_53 b_53 e_53 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_54 c_54 b_54 e_54 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_55 c_55 b_55 e_55 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_56 c_56 b_56 e_56 sub npn13G2v we=0.12u le=2.79u 
Q_pattern_57 c_57 b_57 e_57 sub npn13G2v we=0.12u le=2.79u 
Q_pattern_58 c_58 b_58 e_58 sub npn13G2v we=0.12u le=3.22u 
Q_pattern_59 c_59 b_59 e_59 sub npn13G2v we=0.12u le=3.52u 
Q_pattern_60 c_60 b_60 e_60 sub npn13G2v we=0.12u le=2.55u 
Q_pattern_61 c_61 b_61 e_61 sub npn13G2v we=0.12u le=2.17u 
Q_pattern_62 c_62 b_62 e_62 sub npn13G2v we=0.12u le=4.45u 
Q_pattern_63 c_63 b_63 e_63 sub npn13G2v we=0.12u le=3.14u 
Q_pattern_64 c_64 b_64 e_64 sub npn13G2v we=0.12u le=1.63u 
.ENDS
