*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rppd
Rp1 net1 net2 rppd m=1 l=0.5u w=0.5u
Rp2 net3 net4 rppd m=1 l=1u w=0.5u
Rp3 net5 net6 rppd m=1 l=1.2u w=0.7u
Rp4 net7 net8 rppd m=1 l=1u w=0.5u ps=0.2u b=1
Rp5 net9 net10 rppd m=1 l=1.2u w=0.5u ps=0.2u b=2
.ENDS
