# ------------------------------------------------------
#
#		Copyright 2023 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Thu Jun 12 11:08:54 2025		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_2P_64x32_c2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_2P_64x32_c2 0 0 ;
  SIZE 702.83 BY 74.87 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 425.49 0 425.75 0.26 ;
    END
  END A_DIN[16]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 277.08 0 277.34 0.26 ;
    END
  END A_DIN[15]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 418.35 0 418.61 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 284.22 0 284.48 0.26 ;
    END
  END A_DOUT[15]
  PIN B_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 428.04 0 428.3 0.26 ;
    END
  END B_DIN[16]
  PIN B_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 274.53 0 274.79 0.26 ;
    END
  END B_DIN[15]
  PIN B_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 435.18 0 435.44 0.26 ;
    END
  END B_DOUT[16]
  PIN B_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 267.39 0 267.65 0.26 ;
    END
  END B_DOUT[15]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 683.425 0 687.845 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 665.745 0 670.165 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 648.065 0 652.485 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 630.385 0 634.805 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 612.705 0 617.125 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 595.025 0 599.445 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 577.345 0 581.765 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.665 0 564.085 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 541.985 0 546.405 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 524.305 0 528.725 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.625 0 511.045 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.945 0 493.365 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 471.265 0 475.685 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 453.585 0 458.005 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 435.905 0 440.325 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 418.225 0 422.645 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 388.635 0 391.445 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 378.335 0 381.145 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 362.885 0 365.695 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.585 0 355.395 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.435 0 350.245 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 337.135 0 339.945 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 321.685 0 324.495 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 311.385 0 314.195 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.185 0 284.605 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.505 0 266.925 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 244.825 0 249.245 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 227.145 0 231.565 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 209.465 0 213.885 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 191.785 0 196.205 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.105 0 178.525 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.425 0 160.845 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.745 0 143.165 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 121.065 0 125.485 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 103.385 0 107.805 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.705 0 90.125 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.025 0 72.445 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 50.345 0 54.765 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.665 0 37.085 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 14.985 0 19.405 74.87 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 692.265 0 696.685 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 674.585 0 679.005 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 656.905 0 661.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.225 0 643.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 621.545 0 625.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 603.865 0 608.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.185 0 590.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.505 0 572.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.825 0 555.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.145 0 537.565 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.465 0 519.885 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 497.785 0 502.205 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 480.105 0 484.525 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.425 0 466.845 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 444.745 0 449.165 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.065 0 431.485 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 383.485 0 386.295 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 373.185 0 375.995 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.035 0 370.845 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 357.735 0 360.545 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.285 0 345.095 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 331.985 0 334.795 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.835 0 329.645 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 316.535 0 319.345 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 271.345 0 275.765 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 253.665 0 258.085 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.985 0 240.405 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.305 0 222.725 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.625 0 205.045 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.945 0 187.365 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.265 0 169.685 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.585 0 152.005 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 0 134.325 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 0 116.645 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 0 98.965 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 0 81.285 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 0 63.605 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 0 45.925 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 0 28.245 47.045 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 0 10.565 47.045 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 692.265 53.41 696.685 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 674.585 53.41 679.005 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 656.905 53.41 661.325 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.225 53.41 643.645 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 621.545 53.41 625.965 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 603.865 53.41 608.285 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.185 53.41 590.605 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 568.505 53.41 572.925 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.825 53.41 555.245 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 533.145 53.41 537.565 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.465 53.41 519.885 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 497.785 53.41 502.205 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 480.105 53.41 484.525 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 462.425 53.41 466.845 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 444.745 53.41 449.165 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 427.065 53.41 431.485 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 271.345 53.41 275.765 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 253.665 53.41 258.085 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 235.985 53.41 240.405 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 218.305 53.41 222.725 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.625 53.41 205.045 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.945 53.41 187.365 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 165.265 53.41 169.685 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.585 53.41 152.005 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 129.905 53.41 134.325 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.225 53.41 116.645 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 94.545 53.41 98.965 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.865 53.41 81.285 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.185 53.41 63.605 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 41.505 53.41 45.925 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.825 53.41 28.245 74.87 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.145 53.41 10.565 74.87 ;
    END
  END VDDARRAY!
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 443.17 0 443.43 0.26 ;
    END
  END A_DIN[17]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 259.4 0 259.66 0.26 ;
    END
  END A_DIN[14]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 436.03 0 436.29 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.54 0 266.8 0.26 ;
    END
  END A_DOUT[14]
  PIN B_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 445.72 0 445.98 0.26 ;
    END
  END B_DIN[17]
  PIN B_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 256.85 0 257.11 0.26 ;
    END
  END B_DIN[14]
  PIN B_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 452.86 0 453.12 0.26 ;
    END
  END B_DOUT[17]
  PIN B_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 249.71 0 249.97 0.26 ;
    END
  END B_DOUT[14]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 460.85 0 461.11 0.26 ;
    END
  END A_DIN[18]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 241.72 0 241.98 0.26 ;
    END
  END A_DIN[13]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 453.71 0 453.97 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 248.86 0 249.12 0.26 ;
    END
  END A_DOUT[13]
  PIN B_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 463.4 0 463.66 0.26 ;
    END
  END B_DIN[18]
  PIN B_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 239.17 0 239.43 0.26 ;
    END
  END B_DIN[13]
  PIN B_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 470.54 0 470.8 0.26 ;
    END
  END B_DOUT[18]
  PIN B_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 232.03 0 232.29 0.26 ;
    END
  END B_DOUT[13]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 478.53 0 478.79 0.26 ;
    END
  END A_DIN[19]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 224.04 0 224.3 0.26 ;
    END
  END A_DIN[12]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 471.39 0 471.65 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 231.18 0 231.44 0.26 ;
    END
  END A_DOUT[12]
  PIN B_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 481.08 0 481.34 0.26 ;
    END
  END B_DIN[19]
  PIN B_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221.49 0 221.75 0.26 ;
    END
  END B_DIN[12]
  PIN B_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 488.22 0 488.48 0.26 ;
    END
  END B_DOUT[19]
  PIN B_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 214.35 0 214.61 0.26 ;
    END
  END B_DOUT[12]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 496.21 0 496.47 0.26 ;
    END
  END A_DIN[20]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 206.36 0 206.62 0.26 ;
    END
  END A_DIN[11]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 489.07 0 489.33 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 213.5 0 213.76 0.26 ;
    END
  END A_DOUT[11]
  PIN B_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 498.76 0 499.02 0.26 ;
    END
  END B_DIN[20]
  PIN B_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 203.81 0 204.07 0.26 ;
    END
  END B_DIN[11]
  PIN B_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 505.9 0 506.16 0.26 ;
    END
  END B_DOUT[20]
  PIN B_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 196.67 0 196.93 0.26 ;
    END
  END B_DOUT[11]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 513.89 0 514.15 0.26 ;
    END
  END A_DIN[21]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 188.68 0 188.94 0.26 ;
    END
  END A_DIN[10]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 506.75 0 507.01 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 195.82 0 196.08 0.26 ;
    END
  END A_DOUT[10]
  PIN B_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 516.44 0 516.7 0.26 ;
    END
  END B_DIN[21]
  PIN B_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 186.13 0 186.39 0.26 ;
    END
  END B_DIN[10]
  PIN B_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 523.58 0 523.84 0.26 ;
    END
  END B_DOUT[21]
  PIN B_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.99 0 179.25 0.26 ;
    END
  END B_DOUT[10]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 531.57 0 531.83 0.26 ;
    END
  END A_DIN[22]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 171 0 171.26 0.26 ;
    END
  END A_DIN[9]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 524.43 0 524.69 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 178.14 0 178.4 0.26 ;
    END
  END A_DOUT[9]
  PIN B_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 534.12 0 534.38 0.26 ;
    END
  END B_DIN[22]
  PIN B_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 168.45 0 168.71 0.26 ;
    END
  END B_DIN[9]
  PIN B_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 541.26 0 541.52 0.26 ;
    END
  END B_DOUT[22]
  PIN B_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 161.31 0 161.57 0.26 ;
    END
  END B_DOUT[9]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 549.25 0 549.51 0.26 ;
    END
  END A_DIN[23]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 153.32 0 153.58 0.26 ;
    END
  END A_DIN[8]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 542.11 0 542.37 0.26 ;
    END
  END A_DOUT[23]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 160.46 0 160.72 0.26 ;
    END
  END A_DOUT[8]
  PIN B_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 551.8 0 552.06 0.26 ;
    END
  END B_DIN[23]
  PIN B_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 150.77 0 151.03 0.26 ;
    END
  END B_DIN[8]
  PIN B_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 558.94 0 559.2 0.26 ;
    END
  END B_DOUT[23]
  PIN B_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.63 0 143.89 0.26 ;
    END
  END B_DOUT[8]
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 566.93 0 567.19 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.64 0 135.9 0.26 ;
    END
  END A_DIN[7]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 559.79 0 560.05 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 142.78 0 143.04 0.26 ;
    END
  END A_DOUT[7]
  PIN B_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 569.48 0 569.74 0.26 ;
    END
  END B_DIN[24]
  PIN B_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 133.09 0 133.35 0.26 ;
    END
  END B_DIN[7]
  PIN B_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 576.62 0 576.88 0.26 ;
    END
  END B_DOUT[24]
  PIN B_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.95 0 126.21 0.26 ;
    END
  END B_DOUT[7]
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 584.61 0 584.87 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 117.96 0 118.22 0.26 ;
    END
  END A_DIN[6]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 577.47 0 577.73 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.1 0 125.36 0.26 ;
    END
  END A_DOUT[6]
  PIN B_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 587.16 0 587.42 0.26 ;
    END
  END B_DIN[25]
  PIN B_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 115.41 0 115.67 0.26 ;
    END
  END B_DIN[6]
  PIN B_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 594.3 0 594.56 0.26 ;
    END
  END B_DOUT[25]
  PIN B_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.27 0 108.53 0.26 ;
    END
  END B_DOUT[6]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 602.29 0 602.55 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 100.28 0 100.54 0.26 ;
    END
  END A_DIN[5]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 595.15 0 595.41 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 107.42 0 107.68 0.26 ;
    END
  END A_DOUT[5]
  PIN B_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 604.84 0 605.1 0.26 ;
    END
  END B_DIN[26]
  PIN B_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 97.73 0 97.99 0.26 ;
    END
  END B_DIN[5]
  PIN B_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 611.98 0 612.24 0.26 ;
    END
  END B_DOUT[26]
  PIN B_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 90.59 0 90.85 0.26 ;
    END
  END B_DOUT[5]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 619.97 0 620.23 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.6 0 82.86 0.26 ;
    END
  END A_DIN[4]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 612.83 0 613.09 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.74 0 90 0.26 ;
    END
  END A_DOUT[4]
  PIN B_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 622.52 0 622.78 0.26 ;
    END
  END B_DIN[27]
  PIN B_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 80.05 0 80.31 0.26 ;
    END
  END B_DIN[4]
  PIN B_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 629.66 0 629.92 0.26 ;
    END
  END B_DOUT[27]
  PIN B_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.91 0 73.17 0.26 ;
    END
  END B_DOUT[4]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 637.65 0 637.91 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.92 0 65.18 0.26 ;
    END
  END A_DIN[3]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 630.51 0 630.77 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.06 0 72.32 0.26 ;
    END
  END A_DOUT[3]
  PIN B_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 640.2 0 640.46 0.26 ;
    END
  END B_DIN[28]
  PIN B_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 62.37 0 62.63 0.26 ;
    END
  END B_DIN[3]
  PIN B_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 647.34 0 647.6 0.26 ;
    END
  END B_DOUT[28]
  PIN B_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 55.23 0 55.49 0.26 ;
    END
  END B_DOUT[3]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 655.33 0 655.59 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.24 0 47.5 0.26 ;
    END
  END A_DIN[2]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 648.19 0 648.45 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 54.38 0 54.64 0.26 ;
    END
  END A_DOUT[2]
  PIN B_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 657.88 0 658.14 0.26 ;
    END
  END B_DIN[29]
  PIN B_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.69 0 44.95 0.26 ;
    END
  END B_DIN[2]
  PIN B_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 665.02 0 665.28 0.26 ;
    END
  END B_DOUT[29]
  PIN B_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.55 0 37.81 0.26 ;
    END
  END B_DOUT[2]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 673.01 0 673.27 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 29.56 0 29.82 0.26 ;
    END
  END A_DIN[1]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 665.87 0 666.13 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 36.7 0 36.96 0.26 ;
    END
  END A_DOUT[1]
  PIN B_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 675.56 0 675.82 0.26 ;
    END
  END B_DIN[30]
  PIN B_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 27.01 0 27.27 0.26 ;
    END
  END B_DIN[1]
  PIN B_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 682.7 0 682.96 0.26 ;
    END
  END B_DOUT[30]
  PIN B_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.87 0 20.13 0.26 ;
    END
  END B_DOUT[1]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 690.69 0 690.95 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9091 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.368932 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.88 0 12.14 0.26 ;
    END
  END A_DIN[0]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 683.55 0 683.81 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8256 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 19.02 0 19.28 0.26 ;
    END
  END A_DOUT[0]
  PIN B_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 693.24 0 693.5 0.26 ;
    END
  END B_DIN[31]
  PIN B_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.925 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.469256 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.33 0 9.59 0.26 ;
    END
  END B_DIN[0]
  PIN B_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 700.38 0 700.64 0.26 ;
    END
  END B_DOUT[31]
  PIN B_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.836 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.19 0 2.45 0.26 ;
    END
  END B_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 367.505 0 367.765 0.26 ;
    END
  END A_ADDR[0]
  PIN B_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 335.065 0 335.325 0.26 ;
    END
  END B_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 368.015 0 368.275 0.26 ;
    END
  END A_ADDR[1]
  PIN B_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0851 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 56.097087 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.555 0 334.815 0.26 ;
    END
  END B_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 376.685 0 376.945 0.26 ;
    END
  END A_ADDR[2]
  PIN B_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 325.885 0 326.145 0.26 ;
    END
  END B_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 375.665 0 375.925 0.26 ;
    END
  END A_ADDR[3]
  PIN B_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0819 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.9459 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 21.471247 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 326.905 0 327.165 0.26 ;
    END
  END B_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.285 0 356.545 0.26 ;
    END
  END A_ADDR[4]
  PIN B_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7329 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 74.2589 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 346.285 0 346.545 0.26 ;
    END
  END B_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.265 0 355.525 0.26 ;
    END
  END A_ADDR[5]
  PIN B_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2691 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 66.970874 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 347.305 0 347.565 0.26 ;
    END
  END B_ADDR[5]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 365.975 0 366.235 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 369.545 0 369.805 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 369.035 0 369.295 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 366.485 0 366.745 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 386.885 0 387.145 0.26 ;
    END
  END A_DLY
  PIN B_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 336.595 0 336.855 0.26 ;
    END
  END B_CLK
  PIN B_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.98465 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.745083 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.025 0 333.285 0.26 ;
    END
  END B_REN
  PIN B_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 333.535 0 333.795 0.26 ;
    END
  END B_WEN
  PIN B_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 336.085 0 336.345 0.26 ;
    END
  END B_MEN
  PIN B_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7792 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 23.644788 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 315.685 0 315.945 0.26 ;
    END
  END B_DLY
  OBS
    LAYER Metal1 ;
      RECT 0 0 702.83 74.87 ;
    LAYER Metal2 ;
      RECT 0.31 53.41 0.51 74.84 ;
      RECT 1.135 74.11 1.335 74.84 ;
      RECT 1.545 74.11 1.905 74.84 ;
      RECT 2.115 74.11 2.315 74.84 ;
      RECT 2.19 0.52 2.45 7.78 ;
      RECT 2.7 0.3 2.96 5.235 ;
      RECT 2.77 74.11 2.97 74.84 ;
      RECT 3.21 0 3.47 5.57 ;
      RECT 3.18 74.11 3.54 74.84 ;
      RECT 3.835 74.11 4.035 74.84 ;
      RECT 4.33 74.11 4.69 74.84 ;
      RECT 4.585 0 4.845 6.28 ;
      RECT 4.9 74.11 5.1 74.84 ;
      RECT 5.555 74.11 5.755 74.84 ;
      RECT 5.965 74.11 6.325 74.84 ;
      RECT 6.535 74.11 6.735 74.84 ;
      RECT 6.27 0.18 7.04 0.88 ;
      RECT 7.19 74.11 7.39 74.84 ;
      RECT 7.29 0.3 7.55 8.7 ;
      RECT 7.6 74.11 7.96 74.84 ;
      RECT 8.255 74.11 8.455 74.84 ;
      RECT 8.75 74.11 9.11 74.84 ;
      RECT 9.84 0.155 10.61 0.445 ;
      RECT 9.84 0.155 10.1 8.665 ;
      RECT 10.35 0.155 10.61 8.665 ;
      RECT 9.32 74.11 9.52 74.84 ;
      RECT 9.33 0.52 9.59 9.955 ;
      RECT 9.975 74.11 10.175 74.84 ;
      RECT 10.385 74.11 10.745 74.84 ;
      RECT 10.86 0 11.12 11.315 ;
      RECT 10.955 74.11 11.155 74.84 ;
      RECT 11.37 0 11.63 13.45 ;
      RECT 11.61 74.11 11.81 74.84 ;
      RECT 11.88 0.52 12.14 14.115 ;
      RECT 12.02 74.11 12.38 74.84 ;
      RECT 12.675 74.11 12.875 74.84 ;
      RECT 14.075 0.155 14.845 0.445 ;
      RECT 14.075 0.155 14.335 13.21 ;
      RECT 14.585 0.155 14.845 13.21 ;
      RECT 13.17 74.11 13.53 74.84 ;
      RECT 13.74 74.11 13.94 74.84 ;
      RECT 15.095 0.18 15.865 0.88 ;
      RECT 15.095 0.18 15.355 12.9 ;
      RECT 15.605 0.18 15.865 12.9 ;
      RECT 14.395 74.11 14.595 74.84 ;
      RECT 14.805 74.11 15.165 74.84 ;
      RECT 15.375 74.11 15.575 74.84 ;
      RECT 16.03 74.11 16.23 74.84 ;
      RECT 16.315 0 16.575 2.82 ;
      RECT 16.44 74.11 16.8 74.84 ;
      RECT 17.095 74.11 17.295 74.84 ;
      RECT 17.59 74.11 17.95 74.84 ;
      RECT 17.845 0 18.105 2.82 ;
      RECT 18.16 74.11 18.36 74.84 ;
      RECT 18.815 74.11 19.015 74.84 ;
      RECT 19.02 0.52 19.28 4.315 ;
      RECT 19.225 74.11 19.585 74.84 ;
      RECT 19.795 74.11 19.995 74.84 ;
      RECT 19.87 0.52 20.13 7.78 ;
      RECT 20.38 0.3 20.64 5.235 ;
      RECT 20.45 74.11 20.65 74.84 ;
      RECT 20.89 0 21.15 5.57 ;
      RECT 20.86 74.11 21.22 74.84 ;
      RECT 21.515 74.11 21.715 74.84 ;
      RECT 22.01 74.11 22.37 74.84 ;
      RECT 22.265 0 22.525 6.28 ;
      RECT 22.58 74.11 22.78 74.84 ;
      RECT 23.235 74.11 23.435 74.84 ;
      RECT 23.645 74.11 24.005 74.84 ;
      RECT 24.215 74.11 24.415 74.84 ;
      RECT 23.95 0.18 24.72 0.88 ;
      RECT 24.87 74.11 25.07 74.84 ;
      RECT 24.97 0.3 25.23 8.7 ;
      RECT 25.28 74.11 25.64 74.84 ;
      RECT 25.935 74.11 26.135 74.84 ;
      RECT 26.43 74.11 26.79 74.84 ;
      RECT 27.52 0.155 28.29 0.445 ;
      RECT 27.52 0.155 27.78 8.665 ;
      RECT 28.03 0.155 28.29 8.665 ;
      RECT 27 74.11 27.2 74.84 ;
      RECT 27.01 0.52 27.27 9.955 ;
      RECT 27.655 74.11 27.855 74.84 ;
      RECT 28.065 74.11 28.425 74.84 ;
      RECT 28.54 0 28.8 11.315 ;
      RECT 28.635 74.11 28.835 74.84 ;
      RECT 29.05 0 29.31 13.45 ;
      RECT 29.29 74.11 29.49 74.84 ;
      RECT 29.56 0.52 29.82 14.115 ;
      RECT 29.7 74.11 30.06 74.84 ;
      RECT 30.355 74.11 30.555 74.84 ;
      RECT 31.755 0.155 32.525 0.445 ;
      RECT 31.755 0.155 32.015 13.21 ;
      RECT 32.265 0.155 32.525 13.21 ;
      RECT 30.85 74.11 31.21 74.84 ;
      RECT 31.42 74.11 31.62 74.84 ;
      RECT 32.775 0.18 33.545 0.88 ;
      RECT 32.775 0.18 33.035 12.9 ;
      RECT 33.285 0.18 33.545 12.9 ;
      RECT 32.075 74.11 32.275 74.84 ;
      RECT 32.485 74.11 32.845 74.84 ;
      RECT 33.055 74.11 33.255 74.84 ;
      RECT 33.71 74.11 33.91 74.84 ;
      RECT 33.995 0 34.255 2.82 ;
      RECT 34.12 74.11 34.48 74.84 ;
      RECT 34.775 74.11 34.975 74.84 ;
      RECT 35.27 74.11 35.63 74.84 ;
      RECT 35.525 0 35.785 2.82 ;
      RECT 35.84 74.11 36.04 74.84 ;
      RECT 36.495 74.11 36.695 74.84 ;
      RECT 36.7 0.52 36.96 4.315 ;
      RECT 36.905 74.11 37.265 74.84 ;
      RECT 37.475 74.11 37.675 74.84 ;
      RECT 37.55 0.52 37.81 7.78 ;
      RECT 38.06 0.3 38.32 5.235 ;
      RECT 38.13 74.11 38.33 74.84 ;
      RECT 38.57 0 38.83 5.57 ;
      RECT 38.54 74.11 38.9 74.84 ;
      RECT 39.195 74.11 39.395 74.84 ;
      RECT 39.69 74.11 40.05 74.84 ;
      RECT 39.945 0 40.205 6.28 ;
      RECT 40.26 74.11 40.46 74.84 ;
      RECT 40.915 74.11 41.115 74.84 ;
      RECT 41.325 74.11 41.685 74.84 ;
      RECT 41.895 74.11 42.095 74.84 ;
      RECT 41.63 0.18 42.4 0.88 ;
      RECT 42.55 74.11 42.75 74.84 ;
      RECT 42.65 0.3 42.91 8.7 ;
      RECT 42.96 74.11 43.32 74.84 ;
      RECT 43.615 74.11 43.815 74.84 ;
      RECT 44.11 74.11 44.47 74.84 ;
      RECT 45.2 0.155 45.97 0.445 ;
      RECT 45.2 0.155 45.46 8.665 ;
      RECT 45.71 0.155 45.97 8.665 ;
      RECT 44.68 74.11 44.88 74.84 ;
      RECT 44.69 0.52 44.95 9.955 ;
      RECT 45.335 74.11 45.535 74.84 ;
      RECT 45.745 74.11 46.105 74.84 ;
      RECT 46.22 0 46.48 11.315 ;
      RECT 46.315 74.11 46.515 74.84 ;
      RECT 46.73 0 46.99 13.45 ;
      RECT 46.97 74.11 47.17 74.84 ;
      RECT 47.24 0.52 47.5 14.115 ;
      RECT 47.38 74.11 47.74 74.84 ;
      RECT 48.035 74.11 48.235 74.84 ;
      RECT 49.435 0.155 50.205 0.445 ;
      RECT 49.435 0.155 49.695 13.21 ;
      RECT 49.945 0.155 50.205 13.21 ;
      RECT 48.53 74.11 48.89 74.84 ;
      RECT 49.1 74.11 49.3 74.84 ;
      RECT 50.455 0.18 51.225 0.88 ;
      RECT 50.455 0.18 50.715 12.9 ;
      RECT 50.965 0.18 51.225 12.9 ;
      RECT 49.755 74.11 49.955 74.84 ;
      RECT 50.165 74.11 50.525 74.84 ;
      RECT 50.735 74.11 50.935 74.84 ;
      RECT 51.39 74.11 51.59 74.84 ;
      RECT 51.675 0 51.935 2.82 ;
      RECT 51.8 74.11 52.16 74.84 ;
      RECT 52.455 74.11 52.655 74.84 ;
      RECT 52.95 74.11 53.31 74.84 ;
      RECT 53.205 0 53.465 2.82 ;
      RECT 53.52 74.11 53.72 74.84 ;
      RECT 54.175 74.11 54.375 74.84 ;
      RECT 54.38 0.52 54.64 4.315 ;
      RECT 54.585 74.11 54.945 74.84 ;
      RECT 55.155 74.11 55.355 74.84 ;
      RECT 55.23 0.52 55.49 7.78 ;
      RECT 55.74 0.3 56 5.235 ;
      RECT 55.81 74.11 56.01 74.84 ;
      RECT 56.25 0 56.51 5.57 ;
      RECT 56.22 74.11 56.58 74.84 ;
      RECT 56.875 74.11 57.075 74.84 ;
      RECT 57.37 74.11 57.73 74.84 ;
      RECT 57.625 0 57.885 6.28 ;
      RECT 57.94 74.11 58.14 74.84 ;
      RECT 58.595 74.11 58.795 74.84 ;
      RECT 59.005 74.11 59.365 74.84 ;
      RECT 59.575 74.11 59.775 74.84 ;
      RECT 59.31 0.18 60.08 0.88 ;
      RECT 60.23 74.11 60.43 74.84 ;
      RECT 60.33 0.3 60.59 8.7 ;
      RECT 60.64 74.11 61 74.84 ;
      RECT 61.295 74.11 61.495 74.84 ;
      RECT 61.79 74.11 62.15 74.84 ;
      RECT 62.88 0.155 63.65 0.445 ;
      RECT 62.88 0.155 63.14 8.665 ;
      RECT 63.39 0.155 63.65 8.665 ;
      RECT 62.36 74.11 62.56 74.84 ;
      RECT 62.37 0.52 62.63 9.955 ;
      RECT 63.015 74.11 63.215 74.84 ;
      RECT 63.425 74.11 63.785 74.84 ;
      RECT 63.9 0 64.16 11.315 ;
      RECT 63.995 74.11 64.195 74.84 ;
      RECT 64.41 0 64.67 13.45 ;
      RECT 64.65 74.11 64.85 74.84 ;
      RECT 64.92 0.52 65.18 14.115 ;
      RECT 65.06 74.11 65.42 74.84 ;
      RECT 65.715 74.11 65.915 74.84 ;
      RECT 67.115 0.155 67.885 0.445 ;
      RECT 67.115 0.155 67.375 13.21 ;
      RECT 67.625 0.155 67.885 13.21 ;
      RECT 66.21 74.11 66.57 74.84 ;
      RECT 66.78 74.11 66.98 74.84 ;
      RECT 68.135 0.18 68.905 0.88 ;
      RECT 68.135 0.18 68.395 12.9 ;
      RECT 68.645 0.18 68.905 12.9 ;
      RECT 67.435 74.11 67.635 74.84 ;
      RECT 67.845 74.11 68.205 74.84 ;
      RECT 68.415 74.11 68.615 74.84 ;
      RECT 69.07 74.11 69.27 74.84 ;
      RECT 69.355 0 69.615 2.82 ;
      RECT 69.48 74.11 69.84 74.84 ;
      RECT 70.135 74.11 70.335 74.84 ;
      RECT 70.63 74.11 70.99 74.84 ;
      RECT 70.885 0 71.145 2.82 ;
      RECT 71.2 74.11 71.4 74.84 ;
      RECT 71.855 74.11 72.055 74.84 ;
      RECT 72.06 0.52 72.32 4.315 ;
      RECT 72.265 74.11 72.625 74.84 ;
      RECT 72.835 74.11 73.035 74.84 ;
      RECT 72.91 0.52 73.17 7.78 ;
      RECT 73.42 0.3 73.68 5.235 ;
      RECT 73.49 74.11 73.69 74.84 ;
      RECT 73.93 0 74.19 5.57 ;
      RECT 73.9 74.11 74.26 74.84 ;
      RECT 74.555 74.11 74.755 74.84 ;
      RECT 75.05 74.11 75.41 74.84 ;
      RECT 75.305 0 75.565 6.28 ;
      RECT 75.62 74.11 75.82 74.84 ;
      RECT 76.275 74.11 76.475 74.84 ;
      RECT 76.685 74.11 77.045 74.84 ;
      RECT 77.255 74.11 77.455 74.84 ;
      RECT 76.99 0.18 77.76 0.88 ;
      RECT 77.91 74.11 78.11 74.84 ;
      RECT 78.01 0.3 78.27 8.7 ;
      RECT 78.32 74.11 78.68 74.84 ;
      RECT 78.975 74.11 79.175 74.84 ;
      RECT 79.47 74.11 79.83 74.84 ;
      RECT 80.56 0.155 81.33 0.445 ;
      RECT 80.56 0.155 80.82 8.665 ;
      RECT 81.07 0.155 81.33 8.665 ;
      RECT 80.04 74.11 80.24 74.84 ;
      RECT 80.05 0.52 80.31 9.955 ;
      RECT 80.695 74.11 80.895 74.84 ;
      RECT 81.105 74.11 81.465 74.84 ;
      RECT 81.58 0 81.84 11.315 ;
      RECT 81.675 74.11 81.875 74.84 ;
      RECT 82.09 0 82.35 13.45 ;
      RECT 82.33 74.11 82.53 74.84 ;
      RECT 82.6 0.52 82.86 14.115 ;
      RECT 82.74 74.11 83.1 74.84 ;
      RECT 83.395 74.11 83.595 74.84 ;
      RECT 84.795 0.155 85.565 0.445 ;
      RECT 84.795 0.155 85.055 13.21 ;
      RECT 85.305 0.155 85.565 13.21 ;
      RECT 83.89 74.11 84.25 74.84 ;
      RECT 84.46 74.11 84.66 74.84 ;
      RECT 85.815 0.18 86.585 0.88 ;
      RECT 85.815 0.18 86.075 12.9 ;
      RECT 86.325 0.18 86.585 12.9 ;
      RECT 85.115 74.11 85.315 74.84 ;
      RECT 85.525 74.11 85.885 74.84 ;
      RECT 86.095 74.11 86.295 74.84 ;
      RECT 86.75 74.11 86.95 74.84 ;
      RECT 87.035 0 87.295 2.82 ;
      RECT 87.16 74.11 87.52 74.84 ;
      RECT 87.815 74.11 88.015 74.84 ;
      RECT 88.31 74.11 88.67 74.84 ;
      RECT 88.565 0 88.825 2.82 ;
      RECT 88.88 74.11 89.08 74.84 ;
      RECT 89.535 74.11 89.735 74.84 ;
      RECT 89.74 0.52 90 4.315 ;
      RECT 89.945 74.11 90.305 74.84 ;
      RECT 90.515 74.11 90.715 74.84 ;
      RECT 90.59 0.52 90.85 7.78 ;
      RECT 91.1 0.3 91.36 5.235 ;
      RECT 91.17 74.11 91.37 74.84 ;
      RECT 91.61 0 91.87 5.57 ;
      RECT 91.58 74.11 91.94 74.84 ;
      RECT 92.235 74.11 92.435 74.84 ;
      RECT 92.73 74.11 93.09 74.84 ;
      RECT 92.985 0 93.245 6.28 ;
      RECT 93.3 74.11 93.5 74.84 ;
      RECT 93.955 74.11 94.155 74.84 ;
      RECT 94.365 74.11 94.725 74.84 ;
      RECT 94.935 74.11 95.135 74.84 ;
      RECT 94.67 0.18 95.44 0.88 ;
      RECT 95.59 74.11 95.79 74.84 ;
      RECT 95.69 0.3 95.95 8.7 ;
      RECT 96 74.11 96.36 74.84 ;
      RECT 96.655 74.11 96.855 74.84 ;
      RECT 97.15 74.11 97.51 74.84 ;
      RECT 98.24 0.155 99.01 0.445 ;
      RECT 98.24 0.155 98.5 8.665 ;
      RECT 98.75 0.155 99.01 8.665 ;
      RECT 97.72 74.11 97.92 74.84 ;
      RECT 97.73 0.52 97.99 9.955 ;
      RECT 98.375 74.11 98.575 74.84 ;
      RECT 98.785 74.11 99.145 74.84 ;
      RECT 99.26 0 99.52 11.315 ;
      RECT 99.355 74.11 99.555 74.84 ;
      RECT 99.77 0 100.03 13.45 ;
      RECT 100.01 74.11 100.21 74.84 ;
      RECT 100.28 0.52 100.54 14.115 ;
      RECT 100.42 74.11 100.78 74.84 ;
      RECT 101.075 74.11 101.275 74.84 ;
      RECT 102.475 0.155 103.245 0.445 ;
      RECT 102.475 0.155 102.735 13.21 ;
      RECT 102.985 0.155 103.245 13.21 ;
      RECT 101.57 74.11 101.93 74.84 ;
      RECT 102.14 74.11 102.34 74.84 ;
      RECT 103.495 0.18 104.265 0.88 ;
      RECT 103.495 0.18 103.755 12.9 ;
      RECT 104.005 0.18 104.265 12.9 ;
      RECT 102.795 74.11 102.995 74.84 ;
      RECT 103.205 74.11 103.565 74.84 ;
      RECT 103.775 74.11 103.975 74.84 ;
      RECT 104.43 74.11 104.63 74.84 ;
      RECT 104.715 0 104.975 2.82 ;
      RECT 104.84 74.11 105.2 74.84 ;
      RECT 105.495 74.11 105.695 74.84 ;
      RECT 105.99 74.11 106.35 74.84 ;
      RECT 106.245 0 106.505 2.82 ;
      RECT 106.56 74.11 106.76 74.84 ;
      RECT 107.215 74.11 107.415 74.84 ;
      RECT 107.42 0.52 107.68 4.315 ;
      RECT 107.625 74.11 107.985 74.84 ;
      RECT 108.195 74.11 108.395 74.84 ;
      RECT 108.27 0.52 108.53 7.78 ;
      RECT 108.78 0.3 109.04 5.235 ;
      RECT 108.85 74.11 109.05 74.84 ;
      RECT 109.29 0 109.55 5.57 ;
      RECT 109.26 74.11 109.62 74.84 ;
      RECT 109.915 74.11 110.115 74.84 ;
      RECT 110.41 74.11 110.77 74.84 ;
      RECT 110.665 0 110.925 6.28 ;
      RECT 110.98 74.11 111.18 74.84 ;
      RECT 111.635 74.11 111.835 74.84 ;
      RECT 112.045 74.11 112.405 74.84 ;
      RECT 112.615 74.11 112.815 74.84 ;
      RECT 112.35 0.18 113.12 0.88 ;
      RECT 113.27 74.11 113.47 74.84 ;
      RECT 113.37 0.3 113.63 8.7 ;
      RECT 113.68 74.11 114.04 74.84 ;
      RECT 114.335 74.11 114.535 74.84 ;
      RECT 114.83 74.11 115.19 74.84 ;
      RECT 115.92 0.155 116.69 0.445 ;
      RECT 115.92 0.155 116.18 8.665 ;
      RECT 116.43 0.155 116.69 8.665 ;
      RECT 115.4 74.11 115.6 74.84 ;
      RECT 115.41 0.52 115.67 9.955 ;
      RECT 116.055 74.11 116.255 74.84 ;
      RECT 116.465 74.11 116.825 74.84 ;
      RECT 116.94 0 117.2 11.315 ;
      RECT 117.035 74.11 117.235 74.84 ;
      RECT 117.45 0 117.71 13.45 ;
      RECT 117.69 74.11 117.89 74.84 ;
      RECT 117.96 0.52 118.22 14.115 ;
      RECT 118.1 74.11 118.46 74.84 ;
      RECT 118.755 74.11 118.955 74.84 ;
      RECT 120.155 0.155 120.925 0.445 ;
      RECT 120.155 0.155 120.415 13.21 ;
      RECT 120.665 0.155 120.925 13.21 ;
      RECT 119.25 74.11 119.61 74.84 ;
      RECT 119.82 74.11 120.02 74.84 ;
      RECT 121.175 0.18 121.945 0.88 ;
      RECT 121.175 0.18 121.435 12.9 ;
      RECT 121.685 0.18 121.945 12.9 ;
      RECT 120.475 74.11 120.675 74.84 ;
      RECT 120.885 74.11 121.245 74.84 ;
      RECT 121.455 74.11 121.655 74.84 ;
      RECT 122.11 74.11 122.31 74.84 ;
      RECT 122.395 0 122.655 2.82 ;
      RECT 122.52 74.11 122.88 74.84 ;
      RECT 123.175 74.11 123.375 74.84 ;
      RECT 123.67 74.11 124.03 74.84 ;
      RECT 123.925 0 124.185 2.82 ;
      RECT 124.24 74.11 124.44 74.84 ;
      RECT 124.895 74.11 125.095 74.84 ;
      RECT 125.1 0.52 125.36 4.315 ;
      RECT 125.305 74.11 125.665 74.84 ;
      RECT 125.875 74.11 126.075 74.84 ;
      RECT 125.95 0.52 126.21 7.78 ;
      RECT 126.46 0.3 126.72 5.235 ;
      RECT 126.53 74.11 126.73 74.84 ;
      RECT 126.97 0 127.23 5.57 ;
      RECT 126.94 74.11 127.3 74.84 ;
      RECT 127.595 74.11 127.795 74.84 ;
      RECT 128.09 74.11 128.45 74.84 ;
      RECT 128.345 0 128.605 6.28 ;
      RECT 128.66 74.11 128.86 74.84 ;
      RECT 129.315 74.11 129.515 74.84 ;
      RECT 129.725 74.11 130.085 74.84 ;
      RECT 130.295 74.11 130.495 74.84 ;
      RECT 130.03 0.18 130.8 0.88 ;
      RECT 130.95 74.11 131.15 74.84 ;
      RECT 131.05 0.3 131.31 8.7 ;
      RECT 131.36 74.11 131.72 74.84 ;
      RECT 132.015 74.11 132.215 74.84 ;
      RECT 132.51 74.11 132.87 74.84 ;
      RECT 133.6 0.155 134.37 0.445 ;
      RECT 133.6 0.155 133.86 8.665 ;
      RECT 134.11 0.155 134.37 8.665 ;
      RECT 133.08 74.11 133.28 74.84 ;
      RECT 133.09 0.52 133.35 9.955 ;
      RECT 133.735 74.11 133.935 74.84 ;
      RECT 134.145 74.11 134.505 74.84 ;
      RECT 134.62 0 134.88 11.315 ;
      RECT 134.715 74.11 134.915 74.84 ;
      RECT 135.13 0 135.39 13.45 ;
      RECT 135.37 74.11 135.57 74.84 ;
      RECT 135.64 0.52 135.9 14.115 ;
      RECT 135.78 74.11 136.14 74.84 ;
      RECT 136.435 74.11 136.635 74.84 ;
      RECT 137.835 0.155 138.605 0.445 ;
      RECT 137.835 0.155 138.095 13.21 ;
      RECT 138.345 0.155 138.605 13.21 ;
      RECT 136.93 74.11 137.29 74.84 ;
      RECT 137.5 74.11 137.7 74.84 ;
      RECT 138.855 0.18 139.625 0.88 ;
      RECT 138.855 0.18 139.115 12.9 ;
      RECT 139.365 0.18 139.625 12.9 ;
      RECT 138.155 74.11 138.355 74.84 ;
      RECT 138.565 74.11 138.925 74.84 ;
      RECT 139.135 74.11 139.335 74.84 ;
      RECT 139.79 74.11 139.99 74.84 ;
      RECT 140.075 0 140.335 2.82 ;
      RECT 140.2 74.11 140.56 74.84 ;
      RECT 140.855 74.11 141.055 74.84 ;
      RECT 141.35 74.11 141.71 74.84 ;
      RECT 141.605 0 141.865 2.82 ;
      RECT 141.92 74.11 142.12 74.84 ;
      RECT 142.575 74.11 142.775 74.84 ;
      RECT 142.78 0.52 143.04 4.315 ;
      RECT 142.985 74.11 143.345 74.84 ;
      RECT 143.555 74.11 143.755 74.84 ;
      RECT 143.63 0.52 143.89 7.78 ;
      RECT 144.14 0.3 144.4 5.235 ;
      RECT 144.21 74.11 144.41 74.84 ;
      RECT 144.65 0 144.91 5.57 ;
      RECT 144.62 74.11 144.98 74.84 ;
      RECT 145.275 74.11 145.475 74.84 ;
      RECT 145.77 74.11 146.13 74.84 ;
      RECT 146.025 0 146.285 6.28 ;
      RECT 146.34 74.11 146.54 74.84 ;
      RECT 146.995 74.11 147.195 74.84 ;
      RECT 147.405 74.11 147.765 74.84 ;
      RECT 147.975 74.11 148.175 74.84 ;
      RECT 147.71 0.18 148.48 0.88 ;
      RECT 148.63 74.11 148.83 74.84 ;
      RECT 148.73 0.3 148.99 8.7 ;
      RECT 149.04 74.11 149.4 74.84 ;
      RECT 149.695 74.11 149.895 74.84 ;
      RECT 150.19 74.11 150.55 74.84 ;
      RECT 151.28 0.155 152.05 0.445 ;
      RECT 151.28 0.155 151.54 8.665 ;
      RECT 151.79 0.155 152.05 8.665 ;
      RECT 150.76 74.11 150.96 74.84 ;
      RECT 150.77 0.52 151.03 9.955 ;
      RECT 151.415 74.11 151.615 74.84 ;
      RECT 151.825 74.11 152.185 74.84 ;
      RECT 152.3 0 152.56 11.315 ;
      RECT 152.395 74.11 152.595 74.84 ;
      RECT 152.81 0 153.07 13.45 ;
      RECT 153.05 74.11 153.25 74.84 ;
      RECT 153.32 0.52 153.58 14.115 ;
      RECT 153.46 74.11 153.82 74.84 ;
      RECT 154.115 74.11 154.315 74.84 ;
      RECT 155.515 0.155 156.285 0.445 ;
      RECT 155.515 0.155 155.775 13.21 ;
      RECT 156.025 0.155 156.285 13.21 ;
      RECT 154.61 74.11 154.97 74.84 ;
      RECT 155.18 74.11 155.38 74.84 ;
      RECT 156.535 0.18 157.305 0.88 ;
      RECT 156.535 0.18 156.795 12.9 ;
      RECT 157.045 0.18 157.305 12.9 ;
      RECT 155.835 74.11 156.035 74.84 ;
      RECT 156.245 74.11 156.605 74.84 ;
      RECT 156.815 74.11 157.015 74.84 ;
      RECT 157.47 74.11 157.67 74.84 ;
      RECT 157.755 0 158.015 2.82 ;
      RECT 157.88 74.11 158.24 74.84 ;
      RECT 158.535 74.11 158.735 74.84 ;
      RECT 159.03 74.11 159.39 74.84 ;
      RECT 159.285 0 159.545 2.82 ;
      RECT 159.6 74.11 159.8 74.84 ;
      RECT 160.255 74.11 160.455 74.84 ;
      RECT 160.46 0.52 160.72 4.315 ;
      RECT 160.665 74.11 161.025 74.84 ;
      RECT 161.235 74.11 161.435 74.84 ;
      RECT 161.31 0.52 161.57 7.78 ;
      RECT 161.82 0.3 162.08 5.235 ;
      RECT 161.89 74.11 162.09 74.84 ;
      RECT 162.33 0 162.59 5.57 ;
      RECT 162.3 74.11 162.66 74.84 ;
      RECT 162.955 74.11 163.155 74.84 ;
      RECT 163.45 74.11 163.81 74.84 ;
      RECT 163.705 0 163.965 6.28 ;
      RECT 164.02 74.11 164.22 74.84 ;
      RECT 164.675 74.11 164.875 74.84 ;
      RECT 165.085 74.11 165.445 74.84 ;
      RECT 165.655 74.11 165.855 74.84 ;
      RECT 165.39 0.18 166.16 0.88 ;
      RECT 166.31 74.11 166.51 74.84 ;
      RECT 166.41 0.3 166.67 8.7 ;
      RECT 166.72 74.11 167.08 74.84 ;
      RECT 167.375 74.11 167.575 74.84 ;
      RECT 167.87 74.11 168.23 74.84 ;
      RECT 168.96 0.155 169.73 0.445 ;
      RECT 168.96 0.155 169.22 8.665 ;
      RECT 169.47 0.155 169.73 8.665 ;
      RECT 168.44 74.11 168.64 74.84 ;
      RECT 168.45 0.52 168.71 9.955 ;
      RECT 169.095 74.11 169.295 74.84 ;
      RECT 169.505 74.11 169.865 74.84 ;
      RECT 169.98 0 170.24 11.315 ;
      RECT 170.075 74.11 170.275 74.84 ;
      RECT 170.49 0 170.75 13.45 ;
      RECT 170.73 74.11 170.93 74.84 ;
      RECT 171 0.52 171.26 14.115 ;
      RECT 171.14 74.11 171.5 74.84 ;
      RECT 171.795 74.11 171.995 74.84 ;
      RECT 173.195 0.155 173.965 0.445 ;
      RECT 173.195 0.155 173.455 13.21 ;
      RECT 173.705 0.155 173.965 13.21 ;
      RECT 172.29 74.11 172.65 74.84 ;
      RECT 172.86 74.11 173.06 74.84 ;
      RECT 174.215 0.18 174.985 0.88 ;
      RECT 174.215 0.18 174.475 12.9 ;
      RECT 174.725 0.18 174.985 12.9 ;
      RECT 173.515 74.11 173.715 74.84 ;
      RECT 173.925 74.11 174.285 74.84 ;
      RECT 174.495 74.11 174.695 74.84 ;
      RECT 175.15 74.11 175.35 74.84 ;
      RECT 175.435 0 175.695 2.82 ;
      RECT 175.56 74.11 175.92 74.84 ;
      RECT 176.215 74.11 176.415 74.84 ;
      RECT 176.71 74.11 177.07 74.84 ;
      RECT 176.965 0 177.225 2.82 ;
      RECT 177.28 74.11 177.48 74.84 ;
      RECT 177.935 74.11 178.135 74.84 ;
      RECT 178.14 0.52 178.4 4.315 ;
      RECT 178.345 74.11 178.705 74.84 ;
      RECT 178.915 74.11 179.115 74.84 ;
      RECT 178.99 0.52 179.25 7.78 ;
      RECT 179.5 0.3 179.76 5.235 ;
      RECT 179.57 74.11 179.77 74.84 ;
      RECT 180.01 0 180.27 5.57 ;
      RECT 179.98 74.11 180.34 74.84 ;
      RECT 180.635 74.11 180.835 74.84 ;
      RECT 181.13 74.11 181.49 74.84 ;
      RECT 181.385 0 181.645 6.28 ;
      RECT 181.7 74.11 181.9 74.84 ;
      RECT 182.355 74.11 182.555 74.84 ;
      RECT 182.765 74.11 183.125 74.84 ;
      RECT 183.335 74.11 183.535 74.84 ;
      RECT 183.07 0.18 183.84 0.88 ;
      RECT 183.99 74.11 184.19 74.84 ;
      RECT 184.09 0.3 184.35 8.7 ;
      RECT 184.4 74.11 184.76 74.84 ;
      RECT 185.055 74.11 185.255 74.84 ;
      RECT 185.55 74.11 185.91 74.84 ;
      RECT 186.64 0.155 187.41 0.445 ;
      RECT 186.64 0.155 186.9 8.665 ;
      RECT 187.15 0.155 187.41 8.665 ;
      RECT 186.12 74.11 186.32 74.84 ;
      RECT 186.13 0.52 186.39 9.955 ;
      RECT 186.775 74.11 186.975 74.84 ;
      RECT 187.185 74.11 187.545 74.84 ;
      RECT 187.66 0 187.92 11.315 ;
      RECT 187.755 74.11 187.955 74.84 ;
      RECT 188.17 0 188.43 13.45 ;
      RECT 188.41 74.11 188.61 74.84 ;
      RECT 188.68 0.52 188.94 14.115 ;
      RECT 188.82 74.11 189.18 74.84 ;
      RECT 189.475 74.11 189.675 74.84 ;
      RECT 190.875 0.155 191.645 0.445 ;
      RECT 190.875 0.155 191.135 13.21 ;
      RECT 191.385 0.155 191.645 13.21 ;
      RECT 189.97 74.11 190.33 74.84 ;
      RECT 190.54 74.11 190.74 74.84 ;
      RECT 191.895 0.18 192.665 0.88 ;
      RECT 191.895 0.18 192.155 12.9 ;
      RECT 192.405 0.18 192.665 12.9 ;
      RECT 191.195 74.11 191.395 74.84 ;
      RECT 191.605 74.11 191.965 74.84 ;
      RECT 192.175 74.11 192.375 74.84 ;
      RECT 192.83 74.11 193.03 74.84 ;
      RECT 193.115 0 193.375 2.82 ;
      RECT 193.24 74.11 193.6 74.84 ;
      RECT 193.895 74.11 194.095 74.84 ;
      RECT 194.39 74.11 194.75 74.84 ;
      RECT 194.645 0 194.905 2.82 ;
      RECT 194.96 74.11 195.16 74.84 ;
      RECT 195.615 74.11 195.815 74.84 ;
      RECT 195.82 0.52 196.08 4.315 ;
      RECT 196.025 74.11 196.385 74.84 ;
      RECT 196.595 74.11 196.795 74.84 ;
      RECT 196.67 0.52 196.93 7.78 ;
      RECT 197.18 0.3 197.44 5.235 ;
      RECT 197.25 74.11 197.45 74.84 ;
      RECT 197.69 0 197.95 5.57 ;
      RECT 197.66 74.11 198.02 74.84 ;
      RECT 198.315 74.11 198.515 74.84 ;
      RECT 198.81 74.11 199.17 74.84 ;
      RECT 199.065 0 199.325 6.28 ;
      RECT 199.38 74.11 199.58 74.84 ;
      RECT 200.035 74.11 200.235 74.84 ;
      RECT 200.445 74.11 200.805 74.84 ;
      RECT 201.015 74.11 201.215 74.84 ;
      RECT 200.75 0.18 201.52 0.88 ;
      RECT 201.67 74.11 201.87 74.84 ;
      RECT 201.77 0.3 202.03 8.7 ;
      RECT 202.08 74.11 202.44 74.84 ;
      RECT 202.735 74.11 202.935 74.84 ;
      RECT 203.23 74.11 203.59 74.84 ;
      RECT 204.32 0.155 205.09 0.445 ;
      RECT 204.32 0.155 204.58 8.665 ;
      RECT 204.83 0.155 205.09 8.665 ;
      RECT 203.8 74.11 204 74.84 ;
      RECT 203.81 0.52 204.07 9.955 ;
      RECT 204.455 74.11 204.655 74.84 ;
      RECT 204.865 74.11 205.225 74.84 ;
      RECT 205.34 0 205.6 11.315 ;
      RECT 205.435 74.11 205.635 74.84 ;
      RECT 205.85 0 206.11 13.45 ;
      RECT 206.09 74.11 206.29 74.84 ;
      RECT 206.36 0.52 206.62 14.115 ;
      RECT 206.5 74.11 206.86 74.84 ;
      RECT 207.155 74.11 207.355 74.84 ;
      RECT 208.555 0.155 209.325 0.445 ;
      RECT 208.555 0.155 208.815 13.21 ;
      RECT 209.065 0.155 209.325 13.21 ;
      RECT 207.65 74.11 208.01 74.84 ;
      RECT 208.22 74.11 208.42 74.84 ;
      RECT 209.575 0.18 210.345 0.88 ;
      RECT 209.575 0.18 209.835 12.9 ;
      RECT 210.085 0.18 210.345 12.9 ;
      RECT 208.875 74.11 209.075 74.84 ;
      RECT 209.285 74.11 209.645 74.84 ;
      RECT 209.855 74.11 210.055 74.84 ;
      RECT 210.51 74.11 210.71 74.84 ;
      RECT 210.795 0 211.055 2.82 ;
      RECT 210.92 74.11 211.28 74.84 ;
      RECT 211.575 74.11 211.775 74.84 ;
      RECT 212.07 74.11 212.43 74.84 ;
      RECT 212.325 0 212.585 2.82 ;
      RECT 212.64 74.11 212.84 74.84 ;
      RECT 213.295 74.11 213.495 74.84 ;
      RECT 213.5 0.52 213.76 4.315 ;
      RECT 213.705 74.11 214.065 74.84 ;
      RECT 214.275 74.11 214.475 74.84 ;
      RECT 214.35 0.52 214.61 7.78 ;
      RECT 214.86 0.3 215.12 5.235 ;
      RECT 214.93 74.11 215.13 74.84 ;
      RECT 215.37 0 215.63 5.57 ;
      RECT 215.34 74.11 215.7 74.84 ;
      RECT 215.995 74.11 216.195 74.84 ;
      RECT 216.49 74.11 216.85 74.84 ;
      RECT 216.745 0 217.005 6.28 ;
      RECT 217.06 74.11 217.26 74.84 ;
      RECT 217.715 74.11 217.915 74.84 ;
      RECT 218.125 74.11 218.485 74.84 ;
      RECT 218.695 74.11 218.895 74.84 ;
      RECT 218.43 0.18 219.2 0.88 ;
      RECT 219.35 74.11 219.55 74.84 ;
      RECT 219.45 0.3 219.71 8.7 ;
      RECT 219.76 74.11 220.12 74.84 ;
      RECT 220.415 74.11 220.615 74.84 ;
      RECT 220.91 74.11 221.27 74.84 ;
      RECT 222 0.155 222.77 0.445 ;
      RECT 222 0.155 222.26 8.665 ;
      RECT 222.51 0.155 222.77 8.665 ;
      RECT 221.48 74.11 221.68 74.84 ;
      RECT 221.49 0.52 221.75 9.955 ;
      RECT 222.135 74.11 222.335 74.84 ;
      RECT 222.545 74.11 222.905 74.84 ;
      RECT 223.02 0 223.28 11.315 ;
      RECT 223.115 74.11 223.315 74.84 ;
      RECT 223.53 0 223.79 13.45 ;
      RECT 223.77 74.11 223.97 74.84 ;
      RECT 224.04 0.52 224.3 14.115 ;
      RECT 224.18 74.11 224.54 74.84 ;
      RECT 224.835 74.11 225.035 74.84 ;
      RECT 226.235 0.155 227.005 0.445 ;
      RECT 226.235 0.155 226.495 13.21 ;
      RECT 226.745 0.155 227.005 13.21 ;
      RECT 225.33 74.11 225.69 74.84 ;
      RECT 225.9 74.11 226.1 74.84 ;
      RECT 227.255 0.18 228.025 0.88 ;
      RECT 227.255 0.18 227.515 12.9 ;
      RECT 227.765 0.18 228.025 12.9 ;
      RECT 226.555 74.11 226.755 74.84 ;
      RECT 226.965 74.11 227.325 74.84 ;
      RECT 227.535 74.11 227.735 74.84 ;
      RECT 228.19 74.11 228.39 74.84 ;
      RECT 228.475 0 228.735 2.82 ;
      RECT 228.6 74.11 228.96 74.84 ;
      RECT 229.255 74.11 229.455 74.84 ;
      RECT 229.75 74.11 230.11 74.84 ;
      RECT 230.005 0 230.265 2.82 ;
      RECT 230.32 74.11 230.52 74.84 ;
      RECT 230.975 74.11 231.175 74.84 ;
      RECT 231.18 0.52 231.44 4.315 ;
      RECT 231.385 74.11 231.745 74.84 ;
      RECT 231.955 74.11 232.155 74.84 ;
      RECT 232.03 0.52 232.29 7.78 ;
      RECT 232.54 0.3 232.8 5.235 ;
      RECT 232.61 74.11 232.81 74.84 ;
      RECT 233.05 0 233.31 5.57 ;
      RECT 233.02 74.11 233.38 74.84 ;
      RECT 233.675 74.11 233.875 74.84 ;
      RECT 234.17 74.11 234.53 74.84 ;
      RECT 234.425 0 234.685 6.28 ;
      RECT 234.74 74.11 234.94 74.84 ;
      RECT 235.395 74.11 235.595 74.84 ;
      RECT 235.805 74.11 236.165 74.84 ;
      RECT 236.375 74.11 236.575 74.84 ;
      RECT 236.11 0.18 236.88 0.88 ;
      RECT 237.03 74.11 237.23 74.84 ;
      RECT 237.13 0.3 237.39 8.7 ;
      RECT 237.44 74.11 237.8 74.84 ;
      RECT 238.095 74.11 238.295 74.84 ;
      RECT 238.59 74.11 238.95 74.84 ;
      RECT 239.68 0.155 240.45 0.445 ;
      RECT 239.68 0.155 239.94 8.665 ;
      RECT 240.19 0.155 240.45 8.665 ;
      RECT 239.16 74.11 239.36 74.84 ;
      RECT 239.17 0.52 239.43 9.955 ;
      RECT 239.815 74.11 240.015 74.84 ;
      RECT 240.225 74.11 240.585 74.84 ;
      RECT 240.7 0 240.96 11.315 ;
      RECT 240.795 74.11 240.995 74.84 ;
      RECT 241.21 0 241.47 13.45 ;
      RECT 241.45 74.11 241.65 74.84 ;
      RECT 241.72 0.52 241.98 14.115 ;
      RECT 241.86 74.11 242.22 74.84 ;
      RECT 242.515 74.11 242.715 74.84 ;
      RECT 243.915 0.155 244.685 0.445 ;
      RECT 243.915 0.155 244.175 13.21 ;
      RECT 244.425 0.155 244.685 13.21 ;
      RECT 243.01 74.11 243.37 74.84 ;
      RECT 243.58 74.11 243.78 74.84 ;
      RECT 244.935 0.18 245.705 0.88 ;
      RECT 244.935 0.18 245.195 12.9 ;
      RECT 245.445 0.18 245.705 12.9 ;
      RECT 244.235 74.11 244.435 74.84 ;
      RECT 244.645 74.11 245.005 74.84 ;
      RECT 245.215 74.11 245.415 74.84 ;
      RECT 245.87 74.11 246.07 74.84 ;
      RECT 246.155 0 246.415 2.82 ;
      RECT 246.28 74.11 246.64 74.84 ;
      RECT 246.935 74.11 247.135 74.84 ;
      RECT 247.43 74.11 247.79 74.84 ;
      RECT 247.685 0 247.945 2.82 ;
      RECT 248 74.11 248.2 74.84 ;
      RECT 248.655 74.11 248.855 74.84 ;
      RECT 248.86 0.52 249.12 4.315 ;
      RECT 249.065 74.11 249.425 74.84 ;
      RECT 249.635 74.11 249.835 74.84 ;
      RECT 249.71 0.52 249.97 7.78 ;
      RECT 250.22 0.3 250.48 5.235 ;
      RECT 250.29 74.11 250.49 74.84 ;
      RECT 250.73 0 250.99 5.57 ;
      RECT 250.7 74.11 251.06 74.84 ;
      RECT 251.355 74.11 251.555 74.84 ;
      RECT 251.85 74.11 252.21 74.84 ;
      RECT 252.105 0 252.365 6.28 ;
      RECT 252.42 74.11 252.62 74.84 ;
      RECT 253.075 74.11 253.275 74.84 ;
      RECT 253.485 74.11 253.845 74.84 ;
      RECT 254.055 74.11 254.255 74.84 ;
      RECT 253.79 0.18 254.56 0.88 ;
      RECT 254.71 74.11 254.91 74.84 ;
      RECT 254.81 0.3 255.07 8.7 ;
      RECT 255.12 74.11 255.48 74.84 ;
      RECT 255.775 74.11 255.975 74.84 ;
      RECT 256.27 74.11 256.63 74.84 ;
      RECT 257.36 0.155 258.13 0.445 ;
      RECT 257.36 0.155 257.62 8.665 ;
      RECT 257.87 0.155 258.13 8.665 ;
      RECT 256.84 74.11 257.04 74.84 ;
      RECT 256.85 0.52 257.11 9.955 ;
      RECT 257.495 74.11 257.695 74.84 ;
      RECT 257.905 74.11 258.265 74.84 ;
      RECT 258.38 0 258.64 11.315 ;
      RECT 258.475 74.11 258.675 74.84 ;
      RECT 258.89 0 259.15 13.45 ;
      RECT 259.13 74.11 259.33 74.84 ;
      RECT 259.4 0.52 259.66 14.115 ;
      RECT 259.54 74.11 259.9 74.84 ;
      RECT 260.195 74.11 260.395 74.84 ;
      RECT 261.595 0.155 262.365 0.445 ;
      RECT 261.595 0.155 261.855 13.21 ;
      RECT 262.105 0.155 262.365 13.21 ;
      RECT 260.69 74.11 261.05 74.84 ;
      RECT 261.26 74.11 261.46 74.84 ;
      RECT 262.615 0.18 263.385 0.88 ;
      RECT 262.615 0.18 262.875 12.9 ;
      RECT 263.125 0.18 263.385 12.9 ;
      RECT 261.915 74.11 262.115 74.84 ;
      RECT 262.325 74.11 262.685 74.84 ;
      RECT 262.895 74.11 263.095 74.84 ;
      RECT 263.55 74.11 263.75 74.84 ;
      RECT 263.835 0 264.095 2.82 ;
      RECT 263.96 74.11 264.32 74.84 ;
      RECT 264.615 74.11 264.815 74.84 ;
      RECT 265.11 74.11 265.47 74.84 ;
      RECT 265.365 0 265.625 2.82 ;
      RECT 265.68 74.11 265.88 74.84 ;
      RECT 266.335 74.11 266.535 74.84 ;
      RECT 266.54 0.52 266.8 4.315 ;
      RECT 266.745 74.11 267.105 74.84 ;
      RECT 267.315 74.11 267.515 74.84 ;
      RECT 267.39 0.52 267.65 7.78 ;
      RECT 267.9 0.3 268.16 5.235 ;
      RECT 267.97 74.11 268.17 74.84 ;
      RECT 268.41 0 268.67 5.57 ;
      RECT 268.38 74.11 268.74 74.84 ;
      RECT 269.035 74.11 269.235 74.84 ;
      RECT 269.53 74.11 269.89 74.84 ;
      RECT 269.785 0 270.045 6.28 ;
      RECT 270.1 74.11 270.3 74.84 ;
      RECT 270.755 74.11 270.955 74.84 ;
      RECT 271.165 74.11 271.525 74.84 ;
      RECT 271.735 74.11 271.935 74.84 ;
      RECT 271.47 0.18 272.24 0.88 ;
      RECT 272.39 74.11 272.59 74.84 ;
      RECT 272.49 0.3 272.75 8.7 ;
      RECT 272.8 74.11 273.16 74.84 ;
      RECT 273.455 74.11 273.655 74.84 ;
      RECT 273.95 74.11 274.31 74.84 ;
      RECT 275.04 0.155 275.81 0.445 ;
      RECT 275.04 0.155 275.3 8.665 ;
      RECT 275.55 0.155 275.81 8.665 ;
      RECT 274.52 74.11 274.72 74.84 ;
      RECT 274.53 0.52 274.79 9.955 ;
      RECT 275.175 74.11 275.375 74.84 ;
      RECT 275.585 74.11 275.945 74.84 ;
      RECT 276.06 0 276.32 11.315 ;
      RECT 276.155 74.11 276.355 74.84 ;
      RECT 276.57 0 276.83 13.45 ;
      RECT 276.81 74.11 277.01 74.84 ;
      RECT 277.08 0.52 277.34 14.115 ;
      RECT 277.22 74.11 277.58 74.84 ;
      RECT 277.875 74.11 278.075 74.84 ;
      RECT 279.275 0.155 280.045 0.445 ;
      RECT 279.275 0.155 279.535 13.21 ;
      RECT 279.785 0.155 280.045 13.21 ;
      RECT 278.37 74.11 278.73 74.84 ;
      RECT 278.94 74.11 279.14 74.84 ;
      RECT 280.295 0.18 281.065 0.88 ;
      RECT 280.295 0.18 280.555 12.9 ;
      RECT 280.805 0.18 281.065 12.9 ;
      RECT 279.595 74.11 279.795 74.84 ;
      RECT 280.005 74.11 280.365 74.84 ;
      RECT 280.575 74.11 280.775 74.84 ;
      RECT 281.23 74.11 281.43 74.84 ;
      RECT 281.515 0 281.775 2.82 ;
      RECT 281.64 74.11 282 74.84 ;
      RECT 282.295 74.11 282.495 74.84 ;
      RECT 282.79 74.11 283.15 74.84 ;
      RECT 283.045 0 283.305 2.82 ;
      RECT 283.36 74.11 283.56 74.84 ;
      RECT 284.015 74.11 284.215 74.84 ;
      RECT 284.22 0.52 284.48 4.315 ;
      RECT 285.75 0.17 286.52 0.43 ;
      RECT 285.75 0.17 286.01 8.7 ;
      RECT 286.26 0.17 286.52 8.7 ;
      RECT 286.77 0.18 287.54 0.88 ;
      RECT 286.77 0.18 287.03 8.7 ;
      RECT 287.28 0.18 287.54 8.7 ;
      RECT 287.79 0.17 288.56 0.43 ;
      RECT 287.79 0.17 288.05 8.7 ;
      RECT 288.3 0.17 288.56 8.7 ;
      RECT 288.81 0.18 289.58 0.88 ;
      RECT 288.81 0.18 289.07 8.7 ;
      RECT 289.32 0.18 289.58 8.7 ;
      RECT 289.83 0.17 290.6 0.43 ;
      RECT 289.83 0.17 290.09 8.7 ;
      RECT 290.34 0.17 290.6 8.7 ;
      RECT 290.85 0.18 291.62 0.88 ;
      RECT 290.85 0.18 291.11 8.7 ;
      RECT 291.36 0.18 291.62 8.7 ;
      RECT 291.87 0.17 292.64 0.43 ;
      RECT 291.87 0.17 292.13 8.7 ;
      RECT 292.38 0.17 292.64 8.7 ;
      RECT 292.89 0.18 293.66 0.88 ;
      RECT 292.89 0.18 293.15 8.7 ;
      RECT 293.4 0.18 293.66 8.7 ;
      RECT 293.91 0.17 294.68 0.43 ;
      RECT 293.91 0.17 294.17 8.7 ;
      RECT 294.42 0.17 294.68 8.7 ;
      RECT 294.93 0.18 295.7 0.88 ;
      RECT 294.93 0.18 295.19 8.7 ;
      RECT 295.44 0.18 295.7 8.7 ;
      RECT 295.95 0.17 296.72 0.43 ;
      RECT 295.95 0.17 296.21 8.7 ;
      RECT 296.46 0.17 296.72 8.7 ;
      RECT 296.97 0.18 297.74 0.88 ;
      RECT 296.97 0.18 297.23 8.7 ;
      RECT 297.48 0.18 297.74 8.7 ;
      RECT 297.99 0.17 298.76 0.43 ;
      RECT 297.99 0.17 298.25 8.7 ;
      RECT 298.5 0.17 298.76 8.7 ;
      RECT 299.01 0.18 299.78 0.88 ;
      RECT 299.01 0.18 299.27 8.7 ;
      RECT 299.52 0.18 299.78 8.7 ;
      RECT 300.03 0.17 300.8 0.43 ;
      RECT 300.03 0.17 300.29 8.7 ;
      RECT 300.54 0.17 300.8 8.7 ;
      RECT 301.05 0.18 301.82 0.88 ;
      RECT 301.05 0.18 301.31 8.7 ;
      RECT 301.56 0.18 301.82 8.7 ;
      RECT 302.07 0.17 302.84 0.43 ;
      RECT 302.07 0.17 302.33 8.7 ;
      RECT 302.58 0.17 302.84 8.7 ;
      RECT 303.09 0.18 303.86 0.88 ;
      RECT 303.09 0.18 303.35 8.7 ;
      RECT 303.6 0.18 303.86 8.7 ;
      RECT 304.11 0.17 304.88 0.43 ;
      RECT 304.11 0.17 304.37 8.7 ;
      RECT 304.62 0.17 304.88 8.7 ;
      RECT 305.13 0.18 305.9 0.88 ;
      RECT 305.13 0.18 305.39 8.7 ;
      RECT 305.64 0.18 305.9 8.7 ;
      RECT 306.15 0.17 306.92 0.43 ;
      RECT 306.15 0.17 306.41 8.7 ;
      RECT 306.66 0.17 306.92 8.7 ;
      RECT 307.17 0.18 307.94 0.88 ;
      RECT 307.17 0.18 307.43 8.7 ;
      RECT 307.68 0.18 307.94 8.7 ;
      RECT 308.19 0.17 308.96 0.43 ;
      RECT 308.19 0.17 308.45 8.7 ;
      RECT 308.7 0.17 308.96 8.7 ;
      RECT 309.21 0.18 309.98 0.88 ;
      RECT 309.21 0.18 309.47 8.7 ;
      RECT 309.72 0.18 309.98 8.7 ;
      RECT 284.425 74.11 284.785 74.84 ;
      RECT 284.995 74.11 285.195 74.84 ;
      RECT 311.605 0.18 312.375 0.88 ;
      RECT 311.605 0.18 311.865 8.7 ;
      RECT 312.115 0.18 312.375 8.7 ;
      RECT 312.625 0.17 313.395 0.43 ;
      RECT 312.625 0.17 312.885 8.7 ;
      RECT 313.135 0.17 313.395 8.7 ;
      RECT 285.82 74.03 286.02 74.84 ;
      RECT 310.585 0.3 310.845 8.7 ;
      RECT 314.665 0.18 315.435 0.88 ;
      RECT 314.665 0.18 314.925 8.7 ;
      RECT 315.175 0.18 315.435 8.7 ;
      RECT 311.095 0.3 311.355 8.7 ;
      RECT 313.645 0 313.905 8.7 ;
      RECT 314.155 0 314.415 8.7 ;
      RECT 315.685 0.52 315.945 8.7 ;
      RECT 316.195 0.3 316.455 8.7 ;
      RECT 316.705 0.3 316.965 8.7 ;
      RECT 317.215 0.3 317.475 8.7 ;
      RECT 317.725 0.3 317.985 8.7 ;
      RECT 318.235 0.3 318.495 8.7 ;
      RECT 318.745 0.3 319.005 8.7 ;
      RECT 319.255 0.3 319.515 8.7 ;
      RECT 321.295 0.18 322.065 0.88 ;
      RECT 321.295 0.18 321.555 8.7 ;
      RECT 321.805 0.18 322.065 8.7 ;
      RECT 319.765 0.3 320.025 8.7 ;
      RECT 320.275 0 320.535 8.7 ;
      RECT 320.785 0 321.045 8.7 ;
      RECT 322.315 0 322.575 8.7 ;
      RECT 322.825 0 323.085 8.7 ;
      RECT 323.335 0 323.595 8.7 ;
      RECT 323.845 0 324.105 8.7 ;
      RECT 324.355 0 324.615 8.7 ;
      RECT 324.865 0 325.125 8.7 ;
      RECT 325.375 0 325.635 8.7 ;
      RECT 325.885 0.52 326.145 8.7 ;
      RECT 326.395 0 326.655 8.7 ;
      RECT 326.905 0.52 327.165 8.7 ;
      RECT 327.415 0.3 327.675 8.7 ;
      RECT 327.925 0.3 328.185 8.7 ;
      RECT 328.435 0.3 328.695 8.7 ;
      RECT 328.945 0 329.205 8.7 ;
      RECT 329.455 0 329.715 8.7 ;
      RECT 329.965 0.3 330.225 8.7 ;
      RECT 330.475 0.3 330.735 8.7 ;
      RECT 330.985 0.3 331.245 8.7 ;
      RECT 331.495 0 331.755 8.7 ;
      RECT 332.005 0 332.265 8.7 ;
      RECT 332.515 0.3 332.775 8.7 ;
      RECT 333.025 0.52 333.285 8.7 ;
      RECT 333.535 0.52 333.795 8.7 ;
      RECT 334.045 0 334.305 8.7 ;
      RECT 334.555 0.52 334.815 8.7 ;
      RECT 335.065 0.52 335.325 8.7 ;
      RECT 335.575 0.3 335.835 8.7 ;
      RECT 336.085 0.52 336.345 8.7 ;
      RECT 336.595 0.52 336.855 8.7 ;
      RECT 337.105 0.3 337.365 8.7 ;
      RECT 337.615 0 337.875 8.7 ;
      RECT 339.655 0.17 340.425 0.43 ;
      RECT 339.655 0.17 339.915 8.7 ;
      RECT 340.165 0.17 340.425 8.7 ;
      RECT 338.125 0 338.385 8.7 ;
      RECT 338.635 0.3 338.895 8.7 ;
      RECT 339.145 0.3 339.405 8.7 ;
      RECT 342.205 0.17 342.975 0.43 ;
      RECT 342.205 0.17 342.465 8.7 ;
      RECT 342.715 0.17 342.975 8.7 ;
      RECT 340.675 0.3 340.935 8.7 ;
      RECT 343.735 0.18 344.505 0.88 ;
      RECT 343.735 0.18 343.995 8.7 ;
      RECT 344.245 0.18 344.505 8.7 ;
      RECT 341.185 0.3 341.445 8.7 ;
      RECT 341.695 0.3 341.955 8.7 ;
      RECT 343.225 0.3 343.485 8.7 ;
      RECT 344.755 0 345.015 8.7 ;
      RECT 345.265 0 345.525 8.7 ;
      RECT 345.775 0 346.035 8.7 ;
      RECT 346.285 0.52 346.545 8.7 ;
      RECT 346.795 0 347.055 8.7 ;
      RECT 347.305 0.52 347.565 8.7 ;
      RECT 347.815 0 348.075 8.7 ;
      RECT 348.325 0 348.585 8.7 ;
      RECT 348.835 0.3 349.095 8.7 ;
      RECT 349.345 0.3 349.605 8.7 ;
      RECT 349.855 0 350.115 8.7 ;
      RECT 350.365 0 350.625 8.7 ;
      RECT 350.875 0.3 351.135 8.7 ;
      RECT 351.695 0.3 351.955 8.7 ;
      RECT 352.205 0 352.465 8.7 ;
      RECT 352.715 0 352.975 8.7 ;
      RECT 353.225 0.3 353.485 8.7 ;
      RECT 353.735 0.3 353.995 8.7 ;
      RECT 354.245 0 354.505 8.7 ;
      RECT 354.755 0 355.015 8.7 ;
      RECT 355.265 0.52 355.525 8.7 ;
      RECT 355.775 0 356.035 8.7 ;
      RECT 356.285 0.52 356.545 8.7 ;
      RECT 358.325 0.18 359.095 0.88 ;
      RECT 358.325 0.18 358.585 8.7 ;
      RECT 358.835 0.18 359.095 8.7 ;
      RECT 356.795 0 357.055 8.7 ;
      RECT 359.855 0.17 360.625 0.43 ;
      RECT 359.855 0.17 360.115 8.7 ;
      RECT 360.365 0.17 360.625 8.7 ;
      RECT 357.305 0 357.565 8.7 ;
      RECT 357.815 0 358.075 8.7 ;
      RECT 359.345 0.3 359.605 8.7 ;
      RECT 362.405 0.17 363.175 0.43 ;
      RECT 362.405 0.17 362.665 8.7 ;
      RECT 362.915 0.17 363.175 8.7 ;
      RECT 360.875 0.3 361.135 8.7 ;
      RECT 361.385 0.3 361.645 8.7 ;
      RECT 361.895 0.3 362.155 8.7 ;
      RECT 363.425 0.3 363.685 8.7 ;
      RECT 363.935 0.3 364.195 8.7 ;
      RECT 364.445 0 364.705 8.7 ;
      RECT 364.955 0 365.215 8.7 ;
      RECT 365.465 0.3 365.725 8.7 ;
      RECT 365.975 0.52 366.235 8.7 ;
      RECT 366.485 0.52 366.745 8.7 ;
      RECT 366.995 0.3 367.255 8.7 ;
      RECT 367.505 0.52 367.765 8.7 ;
      RECT 368.015 0.52 368.275 8.7 ;
      RECT 368.525 0 368.785 8.7 ;
      RECT 369.035 0.52 369.295 8.7 ;
      RECT 369.545 0.52 369.805 8.7 ;
      RECT 370.055 0.3 370.315 8.7 ;
      RECT 370.565 0 370.825 8.7 ;
      RECT 371.075 0 371.335 8.7 ;
      RECT 371.585 0.3 371.845 8.7 ;
      RECT 372.095 0.3 372.355 8.7 ;
      RECT 372.605 0.3 372.865 8.7 ;
      RECT 373.115 0 373.375 8.7 ;
      RECT 373.625 0 373.885 8.7 ;
      RECT 374.135 0.3 374.395 8.7 ;
      RECT 374.645 0.3 374.905 8.7 ;
      RECT 375.155 0.3 375.415 8.7 ;
      RECT 375.665 0.52 375.925 8.7 ;
      RECT 376.175 0 376.435 8.7 ;
      RECT 376.685 0.52 376.945 8.7 ;
      RECT 377.195 0 377.455 8.7 ;
      RECT 377.705 0 377.965 8.7 ;
      RECT 378.215 0 378.475 8.7 ;
      RECT 378.725 0 378.985 8.7 ;
      RECT 380.765 0.18 381.535 0.88 ;
      RECT 380.765 0.18 381.025 8.7 ;
      RECT 381.275 0.18 381.535 8.7 ;
      RECT 379.235 0 379.495 8.7 ;
      RECT 379.745 0 380.005 8.7 ;
      RECT 380.255 0 380.515 8.7 ;
      RECT 381.785 0 382.045 8.7 ;
      RECT 382.295 0 382.555 8.7 ;
      RECT 382.805 0.3 383.065 8.7 ;
      RECT 383.315 0.3 383.575 8.7 ;
      RECT 383.825 0.3 384.085 8.7 ;
      RECT 384.335 0.3 384.595 8.7 ;
      RECT 384.845 0.3 385.105 8.7 ;
      RECT 385.355 0.3 385.615 8.7 ;
      RECT 387.395 0.18 388.165 0.88 ;
      RECT 387.395 0.18 387.655 8.7 ;
      RECT 387.905 0.18 388.165 8.7 ;
      RECT 385.865 0.3 386.125 8.7 ;
      RECT 386.375 0.3 386.635 8.7 ;
      RECT 389.435 0.17 390.205 0.43 ;
      RECT 389.435 0.17 389.695 8.7 ;
      RECT 389.945 0.17 390.205 8.7 ;
      RECT 390.455 0.18 391.225 0.88 ;
      RECT 390.455 0.18 390.715 8.7 ;
      RECT 390.965 0.18 391.225 8.7 ;
      RECT 386.885 0.52 387.145 8.7 ;
      RECT 388.415 0 388.675 8.7 ;
      RECT 392.85 0.18 393.62 0.88 ;
      RECT 392.85 0.18 393.11 8.7 ;
      RECT 393.36 0.18 393.62 8.7 ;
      RECT 393.87 0.17 394.64 0.43 ;
      RECT 393.87 0.17 394.13 8.7 ;
      RECT 394.38 0.17 394.64 8.7 ;
      RECT 394.89 0.18 395.66 0.88 ;
      RECT 394.89 0.18 395.15 8.7 ;
      RECT 395.4 0.18 395.66 8.7 ;
      RECT 395.91 0.17 396.68 0.43 ;
      RECT 395.91 0.17 396.17 8.7 ;
      RECT 396.42 0.17 396.68 8.7 ;
      RECT 396.93 0.18 397.7 0.88 ;
      RECT 396.93 0.18 397.19 8.7 ;
      RECT 397.44 0.18 397.7 8.7 ;
      RECT 397.95 0.17 398.72 0.43 ;
      RECT 397.95 0.17 398.21 8.7 ;
      RECT 398.46 0.17 398.72 8.7 ;
      RECT 398.97 0.18 399.74 0.88 ;
      RECT 398.97 0.18 399.23 8.7 ;
      RECT 399.48 0.18 399.74 8.7 ;
      RECT 399.99 0.17 400.76 0.43 ;
      RECT 399.99 0.17 400.25 8.7 ;
      RECT 400.5 0.17 400.76 8.7 ;
      RECT 401.01 0.18 401.78 0.88 ;
      RECT 401.01 0.18 401.27 8.7 ;
      RECT 401.52 0.18 401.78 8.7 ;
      RECT 402.03 0.17 402.8 0.43 ;
      RECT 402.03 0.17 402.29 8.7 ;
      RECT 402.54 0.17 402.8 8.7 ;
      RECT 403.05 0.18 403.82 0.88 ;
      RECT 403.05 0.18 403.31 8.7 ;
      RECT 403.56 0.18 403.82 8.7 ;
      RECT 404.07 0.17 404.84 0.43 ;
      RECT 404.07 0.17 404.33 8.7 ;
      RECT 404.58 0.17 404.84 8.7 ;
      RECT 405.09 0.18 405.86 0.88 ;
      RECT 405.09 0.18 405.35 8.7 ;
      RECT 405.6 0.18 405.86 8.7 ;
      RECT 406.11 0.17 406.88 0.43 ;
      RECT 406.11 0.17 406.37 8.7 ;
      RECT 406.62 0.17 406.88 8.7 ;
      RECT 407.13 0.18 407.9 0.88 ;
      RECT 407.13 0.18 407.39 8.7 ;
      RECT 407.64 0.18 407.9 8.7 ;
      RECT 408.15 0.17 408.92 0.43 ;
      RECT 408.15 0.17 408.41 8.7 ;
      RECT 408.66 0.17 408.92 8.7 ;
      RECT 409.17 0.18 409.94 0.88 ;
      RECT 409.17 0.18 409.43 8.7 ;
      RECT 409.68 0.18 409.94 8.7 ;
      RECT 410.19 0.17 410.96 0.43 ;
      RECT 410.19 0.17 410.45 8.7 ;
      RECT 410.7 0.17 410.96 8.7 ;
      RECT 411.21 0.18 411.98 0.88 ;
      RECT 411.21 0.18 411.47 8.7 ;
      RECT 411.72 0.18 411.98 8.7 ;
      RECT 412.23 0.17 413 0.43 ;
      RECT 412.23 0.17 412.49 8.7 ;
      RECT 412.74 0.17 413 8.7 ;
      RECT 413.25 0.18 414.02 0.88 ;
      RECT 413.25 0.18 413.51 8.7 ;
      RECT 413.76 0.18 414.02 8.7 ;
      RECT 414.27 0.17 415.04 0.43 ;
      RECT 414.27 0.17 414.53 8.7 ;
      RECT 414.78 0.17 415.04 8.7 ;
      RECT 415.29 0.18 416.06 0.88 ;
      RECT 415.29 0.18 415.55 8.7 ;
      RECT 415.8 0.18 416.06 8.7 ;
      RECT 388.925 0 389.185 8.7 ;
      RECT 416.31 0.17 417.08 0.43 ;
      RECT 416.31 0.17 416.57 8.7 ;
      RECT 416.82 0.17 417.08 8.7 ;
      RECT 391.475 0.3 391.735 8.7 ;
      RECT 391.985 0.3 392.245 8.7 ;
      RECT 416.81 74.03 417.01 74.84 ;
      RECT 417.635 74.11 417.835 74.84 ;
      RECT 418.045 74.11 418.405 74.84 ;
      RECT 418.35 0.52 418.61 4.315 ;
      RECT 418.615 74.11 418.815 74.84 ;
      RECT 419.27 74.11 419.47 74.84 ;
      RECT 419.525 0 419.785 2.82 ;
      RECT 419.68 74.11 420.04 74.84 ;
      RECT 420.335 74.11 420.535 74.84 ;
      RECT 420.83 74.11 421.19 74.84 ;
      RECT 421.765 0.18 422.535 0.88 ;
      RECT 421.765 0.18 422.025 12.9 ;
      RECT 422.275 0.18 422.535 12.9 ;
      RECT 421.055 0 421.315 2.82 ;
      RECT 421.4 74.11 421.6 74.84 ;
      RECT 422.785 0.155 423.555 0.445 ;
      RECT 422.785 0.155 423.045 13.21 ;
      RECT 423.295 0.155 423.555 13.21 ;
      RECT 422.055 74.11 422.255 74.84 ;
      RECT 422.465 74.11 422.825 74.84 ;
      RECT 423.035 74.11 423.235 74.84 ;
      RECT 423.69 74.11 423.89 74.84 ;
      RECT 424.1 74.11 424.46 74.84 ;
      RECT 424.755 74.11 424.955 74.84 ;
      RECT 425.25 74.11 425.61 74.84 ;
      RECT 425.49 0.52 425.75 14.115 ;
      RECT 425.82 74.11 426.02 74.84 ;
      RECT 426 0 426.26 13.45 ;
      RECT 426.475 74.11 426.675 74.84 ;
      RECT 427.02 0.155 427.79 0.445 ;
      RECT 427.02 0.155 427.28 8.665 ;
      RECT 427.53 0.155 427.79 8.665 ;
      RECT 426.51 0 426.77 11.315 ;
      RECT 426.885 74.11 427.245 74.84 ;
      RECT 427.455 74.11 427.655 74.84 ;
      RECT 428.04 0.52 428.3 9.955 ;
      RECT 428.11 74.11 428.31 74.84 ;
      RECT 428.52 74.11 428.88 74.84 ;
      RECT 429.175 74.11 429.375 74.84 ;
      RECT 429.67 74.11 430.03 74.84 ;
      RECT 430.08 0.3 430.34 8.7 ;
      RECT 430.24 74.11 430.44 74.84 ;
      RECT 430.895 74.11 431.095 74.84 ;
      RECT 430.59 0.18 431.36 0.88 ;
      RECT 431.305 74.11 431.665 74.84 ;
      RECT 431.875 74.11 432.075 74.84 ;
      RECT 432.53 74.11 432.73 74.84 ;
      RECT 432.785 0 433.045 6.28 ;
      RECT 432.94 74.11 433.3 74.84 ;
      RECT 433.595 74.11 433.795 74.84 ;
      RECT 434.16 0 434.42 5.57 ;
      RECT 434.09 74.11 434.45 74.84 ;
      RECT 434.66 74.11 434.86 74.84 ;
      RECT 434.67 0.3 434.93 5.235 ;
      RECT 435.18 0.52 435.44 7.78 ;
      RECT 435.315 74.11 435.515 74.84 ;
      RECT 435.725 74.11 436.085 74.84 ;
      RECT 436.03 0.52 436.29 4.315 ;
      RECT 436.295 74.11 436.495 74.84 ;
      RECT 436.95 74.11 437.15 74.84 ;
      RECT 437.205 0 437.465 2.82 ;
      RECT 437.36 74.11 437.72 74.84 ;
      RECT 438.015 74.11 438.215 74.84 ;
      RECT 438.51 74.11 438.87 74.84 ;
      RECT 439.445 0.18 440.215 0.88 ;
      RECT 439.445 0.18 439.705 12.9 ;
      RECT 439.955 0.18 440.215 12.9 ;
      RECT 438.735 0 438.995 2.82 ;
      RECT 439.08 74.11 439.28 74.84 ;
      RECT 440.465 0.155 441.235 0.445 ;
      RECT 440.465 0.155 440.725 13.21 ;
      RECT 440.975 0.155 441.235 13.21 ;
      RECT 439.735 74.11 439.935 74.84 ;
      RECT 440.145 74.11 440.505 74.84 ;
      RECT 440.715 74.11 440.915 74.84 ;
      RECT 441.37 74.11 441.57 74.84 ;
      RECT 441.78 74.11 442.14 74.84 ;
      RECT 442.435 74.11 442.635 74.84 ;
      RECT 442.93 74.11 443.29 74.84 ;
      RECT 443.17 0.52 443.43 14.115 ;
      RECT 443.5 74.11 443.7 74.84 ;
      RECT 443.68 0 443.94 13.45 ;
      RECT 444.155 74.11 444.355 74.84 ;
      RECT 444.7 0.155 445.47 0.445 ;
      RECT 444.7 0.155 444.96 8.665 ;
      RECT 445.21 0.155 445.47 8.665 ;
      RECT 444.19 0 444.45 11.315 ;
      RECT 444.565 74.11 444.925 74.84 ;
      RECT 445.135 74.11 445.335 74.84 ;
      RECT 445.72 0.52 445.98 9.955 ;
      RECT 445.79 74.11 445.99 74.84 ;
      RECT 446.2 74.11 446.56 74.84 ;
      RECT 446.855 74.11 447.055 74.84 ;
      RECT 447.35 74.11 447.71 74.84 ;
      RECT 447.76 0.3 448.02 8.7 ;
      RECT 447.92 74.11 448.12 74.84 ;
      RECT 448.575 74.11 448.775 74.84 ;
      RECT 448.27 0.18 449.04 0.88 ;
      RECT 448.985 74.11 449.345 74.84 ;
      RECT 449.555 74.11 449.755 74.84 ;
      RECT 450.21 74.11 450.41 74.84 ;
      RECT 450.465 0 450.725 6.28 ;
      RECT 450.62 74.11 450.98 74.84 ;
      RECT 451.275 74.11 451.475 74.84 ;
      RECT 451.84 0 452.1 5.57 ;
      RECT 451.77 74.11 452.13 74.84 ;
      RECT 452.34 74.11 452.54 74.84 ;
      RECT 452.35 0.3 452.61 5.235 ;
      RECT 452.86 0.52 453.12 7.78 ;
      RECT 452.995 74.11 453.195 74.84 ;
      RECT 453.405 74.11 453.765 74.84 ;
      RECT 453.71 0.52 453.97 4.315 ;
      RECT 453.975 74.11 454.175 74.84 ;
      RECT 454.63 74.11 454.83 74.84 ;
      RECT 454.885 0 455.145 2.82 ;
      RECT 455.04 74.11 455.4 74.84 ;
      RECT 455.695 74.11 455.895 74.84 ;
      RECT 456.19 74.11 456.55 74.84 ;
      RECT 457.125 0.18 457.895 0.88 ;
      RECT 457.125 0.18 457.385 12.9 ;
      RECT 457.635 0.18 457.895 12.9 ;
      RECT 456.415 0 456.675 2.82 ;
      RECT 456.76 74.11 456.96 74.84 ;
      RECT 458.145 0.155 458.915 0.445 ;
      RECT 458.145 0.155 458.405 13.21 ;
      RECT 458.655 0.155 458.915 13.21 ;
      RECT 457.415 74.11 457.615 74.84 ;
      RECT 457.825 74.11 458.185 74.84 ;
      RECT 458.395 74.11 458.595 74.84 ;
      RECT 459.05 74.11 459.25 74.84 ;
      RECT 459.46 74.11 459.82 74.84 ;
      RECT 460.115 74.11 460.315 74.84 ;
      RECT 460.61 74.11 460.97 74.84 ;
      RECT 460.85 0.52 461.11 14.115 ;
      RECT 461.18 74.11 461.38 74.84 ;
      RECT 461.36 0 461.62 13.45 ;
      RECT 461.835 74.11 462.035 74.84 ;
      RECT 462.38 0.155 463.15 0.445 ;
      RECT 462.38 0.155 462.64 8.665 ;
      RECT 462.89 0.155 463.15 8.665 ;
      RECT 461.87 0 462.13 11.315 ;
      RECT 462.245 74.11 462.605 74.84 ;
      RECT 462.815 74.11 463.015 74.84 ;
      RECT 463.4 0.52 463.66 9.955 ;
      RECT 463.47 74.11 463.67 74.84 ;
      RECT 463.88 74.11 464.24 74.84 ;
      RECT 464.535 74.11 464.735 74.84 ;
      RECT 465.03 74.11 465.39 74.84 ;
      RECT 465.44 0.3 465.7 8.7 ;
      RECT 465.6 74.11 465.8 74.84 ;
      RECT 466.255 74.11 466.455 74.84 ;
      RECT 465.95 0.18 466.72 0.88 ;
      RECT 466.665 74.11 467.025 74.84 ;
      RECT 467.235 74.11 467.435 74.84 ;
      RECT 467.89 74.11 468.09 74.84 ;
      RECT 468.145 0 468.405 6.28 ;
      RECT 468.3 74.11 468.66 74.84 ;
      RECT 468.955 74.11 469.155 74.84 ;
      RECT 469.52 0 469.78 5.57 ;
      RECT 469.45 74.11 469.81 74.84 ;
      RECT 470.02 74.11 470.22 74.84 ;
      RECT 470.03 0.3 470.29 5.235 ;
      RECT 470.54 0.52 470.8 7.78 ;
      RECT 470.675 74.11 470.875 74.84 ;
      RECT 471.085 74.11 471.445 74.84 ;
      RECT 471.39 0.52 471.65 4.315 ;
      RECT 471.655 74.11 471.855 74.84 ;
      RECT 472.31 74.11 472.51 74.84 ;
      RECT 472.565 0 472.825 2.82 ;
      RECT 472.72 74.11 473.08 74.84 ;
      RECT 473.375 74.11 473.575 74.84 ;
      RECT 473.87 74.11 474.23 74.84 ;
      RECT 474.805 0.18 475.575 0.88 ;
      RECT 474.805 0.18 475.065 12.9 ;
      RECT 475.315 0.18 475.575 12.9 ;
      RECT 474.095 0 474.355 2.82 ;
      RECT 474.44 74.11 474.64 74.84 ;
      RECT 475.825 0.155 476.595 0.445 ;
      RECT 475.825 0.155 476.085 13.21 ;
      RECT 476.335 0.155 476.595 13.21 ;
      RECT 475.095 74.11 475.295 74.84 ;
      RECT 475.505 74.11 475.865 74.84 ;
      RECT 476.075 74.11 476.275 74.84 ;
      RECT 476.73 74.11 476.93 74.84 ;
      RECT 477.14 74.11 477.5 74.84 ;
      RECT 477.795 74.11 477.995 74.84 ;
      RECT 478.29 74.11 478.65 74.84 ;
      RECT 478.53 0.52 478.79 14.115 ;
      RECT 478.86 74.11 479.06 74.84 ;
      RECT 479.04 0 479.3 13.45 ;
      RECT 479.515 74.11 479.715 74.84 ;
      RECT 480.06 0.155 480.83 0.445 ;
      RECT 480.06 0.155 480.32 8.665 ;
      RECT 480.57 0.155 480.83 8.665 ;
      RECT 479.55 0 479.81 11.315 ;
      RECT 479.925 74.11 480.285 74.84 ;
      RECT 480.495 74.11 480.695 74.84 ;
      RECT 481.08 0.52 481.34 9.955 ;
      RECT 481.15 74.11 481.35 74.84 ;
      RECT 481.56 74.11 481.92 74.84 ;
      RECT 482.215 74.11 482.415 74.84 ;
      RECT 482.71 74.11 483.07 74.84 ;
      RECT 483.12 0.3 483.38 8.7 ;
      RECT 483.28 74.11 483.48 74.84 ;
      RECT 483.935 74.11 484.135 74.84 ;
      RECT 483.63 0.18 484.4 0.88 ;
      RECT 484.345 74.11 484.705 74.84 ;
      RECT 484.915 74.11 485.115 74.84 ;
      RECT 485.57 74.11 485.77 74.84 ;
      RECT 485.825 0 486.085 6.28 ;
      RECT 485.98 74.11 486.34 74.84 ;
      RECT 486.635 74.11 486.835 74.84 ;
      RECT 487.2 0 487.46 5.57 ;
      RECT 487.13 74.11 487.49 74.84 ;
      RECT 487.7 74.11 487.9 74.84 ;
      RECT 487.71 0.3 487.97 5.235 ;
      RECT 488.22 0.52 488.48 7.78 ;
      RECT 488.355 74.11 488.555 74.84 ;
      RECT 488.765 74.11 489.125 74.84 ;
      RECT 489.07 0.52 489.33 4.315 ;
      RECT 489.335 74.11 489.535 74.84 ;
      RECT 489.99 74.11 490.19 74.84 ;
      RECT 490.245 0 490.505 2.82 ;
      RECT 490.4 74.11 490.76 74.84 ;
      RECT 491.055 74.11 491.255 74.84 ;
      RECT 491.55 74.11 491.91 74.84 ;
      RECT 492.485 0.18 493.255 0.88 ;
      RECT 492.485 0.18 492.745 12.9 ;
      RECT 492.995 0.18 493.255 12.9 ;
      RECT 491.775 0 492.035 2.82 ;
      RECT 492.12 74.11 492.32 74.84 ;
      RECT 493.505 0.155 494.275 0.445 ;
      RECT 493.505 0.155 493.765 13.21 ;
      RECT 494.015 0.155 494.275 13.21 ;
      RECT 492.775 74.11 492.975 74.84 ;
      RECT 493.185 74.11 493.545 74.84 ;
      RECT 493.755 74.11 493.955 74.84 ;
      RECT 494.41 74.11 494.61 74.84 ;
      RECT 494.82 74.11 495.18 74.84 ;
      RECT 495.475 74.11 495.675 74.84 ;
      RECT 495.97 74.11 496.33 74.84 ;
      RECT 496.21 0.52 496.47 14.115 ;
      RECT 496.54 74.11 496.74 74.84 ;
      RECT 496.72 0 496.98 13.45 ;
      RECT 497.195 74.11 497.395 74.84 ;
      RECT 497.74 0.155 498.51 0.445 ;
      RECT 497.74 0.155 498 8.665 ;
      RECT 498.25 0.155 498.51 8.665 ;
      RECT 497.23 0 497.49 11.315 ;
      RECT 497.605 74.11 497.965 74.84 ;
      RECT 498.175 74.11 498.375 74.84 ;
      RECT 498.76 0.52 499.02 9.955 ;
      RECT 498.83 74.11 499.03 74.84 ;
      RECT 499.24 74.11 499.6 74.84 ;
      RECT 499.895 74.11 500.095 74.84 ;
      RECT 500.39 74.11 500.75 74.84 ;
      RECT 500.8 0.3 501.06 8.7 ;
      RECT 500.96 74.11 501.16 74.84 ;
      RECT 501.615 74.11 501.815 74.84 ;
      RECT 501.31 0.18 502.08 0.88 ;
      RECT 502.025 74.11 502.385 74.84 ;
      RECT 502.595 74.11 502.795 74.84 ;
      RECT 503.25 74.11 503.45 74.84 ;
      RECT 503.505 0 503.765 6.28 ;
      RECT 503.66 74.11 504.02 74.84 ;
      RECT 504.315 74.11 504.515 74.84 ;
      RECT 504.88 0 505.14 5.57 ;
      RECT 504.81 74.11 505.17 74.84 ;
      RECT 505.38 74.11 505.58 74.84 ;
      RECT 505.39 0.3 505.65 5.235 ;
      RECT 505.9 0.52 506.16 7.78 ;
      RECT 506.035 74.11 506.235 74.84 ;
      RECT 506.445 74.11 506.805 74.84 ;
      RECT 506.75 0.52 507.01 4.315 ;
      RECT 507.015 74.11 507.215 74.84 ;
      RECT 507.67 74.11 507.87 74.84 ;
      RECT 507.925 0 508.185 2.82 ;
      RECT 508.08 74.11 508.44 74.84 ;
      RECT 508.735 74.11 508.935 74.84 ;
      RECT 509.23 74.11 509.59 74.84 ;
      RECT 510.165 0.18 510.935 0.88 ;
      RECT 510.165 0.18 510.425 12.9 ;
      RECT 510.675 0.18 510.935 12.9 ;
      RECT 509.455 0 509.715 2.82 ;
      RECT 509.8 74.11 510 74.84 ;
      RECT 511.185 0.155 511.955 0.445 ;
      RECT 511.185 0.155 511.445 13.21 ;
      RECT 511.695 0.155 511.955 13.21 ;
      RECT 510.455 74.11 510.655 74.84 ;
      RECT 510.865 74.11 511.225 74.84 ;
      RECT 511.435 74.11 511.635 74.84 ;
      RECT 512.09 74.11 512.29 74.84 ;
      RECT 512.5 74.11 512.86 74.84 ;
      RECT 513.155 74.11 513.355 74.84 ;
      RECT 513.65 74.11 514.01 74.84 ;
      RECT 513.89 0.52 514.15 14.115 ;
      RECT 514.22 74.11 514.42 74.84 ;
      RECT 514.4 0 514.66 13.45 ;
      RECT 514.875 74.11 515.075 74.84 ;
      RECT 515.42 0.155 516.19 0.445 ;
      RECT 515.42 0.155 515.68 8.665 ;
      RECT 515.93 0.155 516.19 8.665 ;
      RECT 514.91 0 515.17 11.315 ;
      RECT 515.285 74.11 515.645 74.84 ;
      RECT 515.855 74.11 516.055 74.84 ;
      RECT 516.44 0.52 516.7 9.955 ;
      RECT 516.51 74.11 516.71 74.84 ;
      RECT 516.92 74.11 517.28 74.84 ;
      RECT 517.575 74.11 517.775 74.84 ;
      RECT 518.07 74.11 518.43 74.84 ;
      RECT 518.48 0.3 518.74 8.7 ;
      RECT 518.64 74.11 518.84 74.84 ;
      RECT 519.295 74.11 519.495 74.84 ;
      RECT 518.99 0.18 519.76 0.88 ;
      RECT 519.705 74.11 520.065 74.84 ;
      RECT 520.275 74.11 520.475 74.84 ;
      RECT 520.93 74.11 521.13 74.84 ;
      RECT 521.185 0 521.445 6.28 ;
      RECT 521.34 74.11 521.7 74.84 ;
      RECT 521.995 74.11 522.195 74.84 ;
      RECT 522.56 0 522.82 5.57 ;
      RECT 522.49 74.11 522.85 74.84 ;
      RECT 523.06 74.11 523.26 74.84 ;
      RECT 523.07 0.3 523.33 5.235 ;
      RECT 523.58 0.52 523.84 7.78 ;
      RECT 523.715 74.11 523.915 74.84 ;
      RECT 524.125 74.11 524.485 74.84 ;
      RECT 524.43 0.52 524.69 4.315 ;
      RECT 524.695 74.11 524.895 74.84 ;
      RECT 525.35 74.11 525.55 74.84 ;
      RECT 525.605 0 525.865 2.82 ;
      RECT 525.76 74.11 526.12 74.84 ;
      RECT 526.415 74.11 526.615 74.84 ;
      RECT 526.91 74.11 527.27 74.84 ;
      RECT 527.845 0.18 528.615 0.88 ;
      RECT 527.845 0.18 528.105 12.9 ;
      RECT 528.355 0.18 528.615 12.9 ;
      RECT 527.135 0 527.395 2.82 ;
      RECT 527.48 74.11 527.68 74.84 ;
      RECT 528.865 0.155 529.635 0.445 ;
      RECT 528.865 0.155 529.125 13.21 ;
      RECT 529.375 0.155 529.635 13.21 ;
      RECT 528.135 74.11 528.335 74.84 ;
      RECT 528.545 74.11 528.905 74.84 ;
      RECT 529.115 74.11 529.315 74.84 ;
      RECT 529.77 74.11 529.97 74.84 ;
      RECT 530.18 74.11 530.54 74.84 ;
      RECT 530.835 74.11 531.035 74.84 ;
      RECT 531.33 74.11 531.69 74.84 ;
      RECT 531.57 0.52 531.83 14.115 ;
      RECT 531.9 74.11 532.1 74.84 ;
      RECT 532.08 0 532.34 13.45 ;
      RECT 532.555 74.11 532.755 74.84 ;
      RECT 533.1 0.155 533.87 0.445 ;
      RECT 533.1 0.155 533.36 8.665 ;
      RECT 533.61 0.155 533.87 8.665 ;
      RECT 532.59 0 532.85 11.315 ;
      RECT 532.965 74.11 533.325 74.84 ;
      RECT 533.535 74.11 533.735 74.84 ;
      RECT 534.12 0.52 534.38 9.955 ;
      RECT 534.19 74.11 534.39 74.84 ;
      RECT 534.6 74.11 534.96 74.84 ;
      RECT 535.255 74.11 535.455 74.84 ;
      RECT 535.75 74.11 536.11 74.84 ;
      RECT 536.16 0.3 536.42 8.7 ;
      RECT 536.32 74.11 536.52 74.84 ;
      RECT 536.975 74.11 537.175 74.84 ;
      RECT 536.67 0.18 537.44 0.88 ;
      RECT 537.385 74.11 537.745 74.84 ;
      RECT 537.955 74.11 538.155 74.84 ;
      RECT 538.61 74.11 538.81 74.84 ;
      RECT 538.865 0 539.125 6.28 ;
      RECT 539.02 74.11 539.38 74.84 ;
      RECT 539.675 74.11 539.875 74.84 ;
      RECT 540.24 0 540.5 5.57 ;
      RECT 540.17 74.11 540.53 74.84 ;
      RECT 540.74 74.11 540.94 74.84 ;
      RECT 540.75 0.3 541.01 5.235 ;
      RECT 541.26 0.52 541.52 7.78 ;
      RECT 541.395 74.11 541.595 74.84 ;
      RECT 541.805 74.11 542.165 74.84 ;
      RECT 542.11 0.52 542.37 4.315 ;
      RECT 542.375 74.11 542.575 74.84 ;
      RECT 543.03 74.11 543.23 74.84 ;
      RECT 543.285 0 543.545 2.82 ;
      RECT 543.44 74.11 543.8 74.84 ;
      RECT 544.095 74.11 544.295 74.84 ;
      RECT 544.59 74.11 544.95 74.84 ;
      RECT 545.525 0.18 546.295 0.88 ;
      RECT 545.525 0.18 545.785 12.9 ;
      RECT 546.035 0.18 546.295 12.9 ;
      RECT 544.815 0 545.075 2.82 ;
      RECT 545.16 74.11 545.36 74.84 ;
      RECT 546.545 0.155 547.315 0.445 ;
      RECT 546.545 0.155 546.805 13.21 ;
      RECT 547.055 0.155 547.315 13.21 ;
      RECT 545.815 74.11 546.015 74.84 ;
      RECT 546.225 74.11 546.585 74.84 ;
      RECT 546.795 74.11 546.995 74.84 ;
      RECT 547.45 74.11 547.65 74.84 ;
      RECT 547.86 74.11 548.22 74.84 ;
      RECT 548.515 74.11 548.715 74.84 ;
      RECT 549.01 74.11 549.37 74.84 ;
      RECT 549.25 0.52 549.51 14.115 ;
      RECT 549.58 74.11 549.78 74.84 ;
      RECT 549.76 0 550.02 13.45 ;
      RECT 550.235 74.11 550.435 74.84 ;
      RECT 550.78 0.155 551.55 0.445 ;
      RECT 550.78 0.155 551.04 8.665 ;
      RECT 551.29 0.155 551.55 8.665 ;
      RECT 550.27 0 550.53 11.315 ;
      RECT 550.645 74.11 551.005 74.84 ;
      RECT 551.215 74.11 551.415 74.84 ;
      RECT 551.8 0.52 552.06 9.955 ;
      RECT 551.87 74.11 552.07 74.84 ;
      RECT 552.28 74.11 552.64 74.84 ;
      RECT 552.935 74.11 553.135 74.84 ;
      RECT 553.43 74.11 553.79 74.84 ;
      RECT 553.84 0.3 554.1 8.7 ;
      RECT 554 74.11 554.2 74.84 ;
      RECT 554.655 74.11 554.855 74.84 ;
      RECT 554.35 0.18 555.12 0.88 ;
      RECT 555.065 74.11 555.425 74.84 ;
      RECT 555.635 74.11 555.835 74.84 ;
      RECT 556.29 74.11 556.49 74.84 ;
      RECT 556.545 0 556.805 6.28 ;
      RECT 556.7 74.11 557.06 74.84 ;
      RECT 557.355 74.11 557.555 74.84 ;
      RECT 557.92 0 558.18 5.57 ;
      RECT 557.85 74.11 558.21 74.84 ;
      RECT 558.42 74.11 558.62 74.84 ;
      RECT 558.43 0.3 558.69 5.235 ;
      RECT 558.94 0.52 559.2 7.78 ;
      RECT 559.075 74.11 559.275 74.84 ;
      RECT 559.485 74.11 559.845 74.84 ;
      RECT 559.79 0.52 560.05 4.315 ;
      RECT 560.055 74.11 560.255 74.84 ;
      RECT 560.71 74.11 560.91 74.84 ;
      RECT 560.965 0 561.225 2.82 ;
      RECT 561.12 74.11 561.48 74.84 ;
      RECT 561.775 74.11 561.975 74.84 ;
      RECT 562.27 74.11 562.63 74.84 ;
      RECT 563.205 0.18 563.975 0.88 ;
      RECT 563.205 0.18 563.465 12.9 ;
      RECT 563.715 0.18 563.975 12.9 ;
      RECT 562.495 0 562.755 2.82 ;
      RECT 562.84 74.11 563.04 74.84 ;
      RECT 564.225 0.155 564.995 0.445 ;
      RECT 564.225 0.155 564.485 13.21 ;
      RECT 564.735 0.155 564.995 13.21 ;
      RECT 563.495 74.11 563.695 74.84 ;
      RECT 563.905 74.11 564.265 74.84 ;
      RECT 564.475 74.11 564.675 74.84 ;
      RECT 565.13 74.11 565.33 74.84 ;
      RECT 565.54 74.11 565.9 74.84 ;
      RECT 566.195 74.11 566.395 74.84 ;
      RECT 566.69 74.11 567.05 74.84 ;
      RECT 566.93 0.52 567.19 14.115 ;
      RECT 567.26 74.11 567.46 74.84 ;
      RECT 567.44 0 567.7 13.45 ;
      RECT 567.915 74.11 568.115 74.84 ;
      RECT 568.46 0.155 569.23 0.445 ;
      RECT 568.46 0.155 568.72 8.665 ;
      RECT 568.97 0.155 569.23 8.665 ;
      RECT 567.95 0 568.21 11.315 ;
      RECT 568.325 74.11 568.685 74.84 ;
      RECT 568.895 74.11 569.095 74.84 ;
      RECT 569.48 0.52 569.74 9.955 ;
      RECT 569.55 74.11 569.75 74.84 ;
      RECT 569.96 74.11 570.32 74.84 ;
      RECT 570.615 74.11 570.815 74.84 ;
      RECT 571.11 74.11 571.47 74.84 ;
      RECT 571.52 0.3 571.78 8.7 ;
      RECT 571.68 74.11 571.88 74.84 ;
      RECT 572.335 74.11 572.535 74.84 ;
      RECT 572.03 0.18 572.8 0.88 ;
      RECT 572.745 74.11 573.105 74.84 ;
      RECT 573.315 74.11 573.515 74.84 ;
      RECT 573.97 74.11 574.17 74.84 ;
      RECT 574.225 0 574.485 6.28 ;
      RECT 574.38 74.11 574.74 74.84 ;
      RECT 575.035 74.11 575.235 74.84 ;
      RECT 575.6 0 575.86 5.57 ;
      RECT 575.53 74.11 575.89 74.84 ;
      RECT 576.1 74.11 576.3 74.84 ;
      RECT 576.11 0.3 576.37 5.235 ;
      RECT 576.62 0.52 576.88 7.78 ;
      RECT 576.755 74.11 576.955 74.84 ;
      RECT 577.165 74.11 577.525 74.84 ;
      RECT 577.47 0.52 577.73 4.315 ;
      RECT 577.735 74.11 577.935 74.84 ;
      RECT 578.39 74.11 578.59 74.84 ;
      RECT 578.645 0 578.905 2.82 ;
      RECT 578.8 74.11 579.16 74.84 ;
      RECT 579.455 74.11 579.655 74.84 ;
      RECT 579.95 74.11 580.31 74.84 ;
      RECT 580.885 0.18 581.655 0.88 ;
      RECT 580.885 0.18 581.145 12.9 ;
      RECT 581.395 0.18 581.655 12.9 ;
      RECT 580.175 0 580.435 2.82 ;
      RECT 580.52 74.11 580.72 74.84 ;
      RECT 581.905 0.155 582.675 0.445 ;
      RECT 581.905 0.155 582.165 13.21 ;
      RECT 582.415 0.155 582.675 13.21 ;
      RECT 581.175 74.11 581.375 74.84 ;
      RECT 581.585 74.11 581.945 74.84 ;
      RECT 582.155 74.11 582.355 74.84 ;
      RECT 582.81 74.11 583.01 74.84 ;
      RECT 583.22 74.11 583.58 74.84 ;
      RECT 583.875 74.11 584.075 74.84 ;
      RECT 584.37 74.11 584.73 74.84 ;
      RECT 584.61 0.52 584.87 14.115 ;
      RECT 584.94 74.11 585.14 74.84 ;
      RECT 585.12 0 585.38 13.45 ;
      RECT 585.595 74.11 585.795 74.84 ;
      RECT 586.14 0.155 586.91 0.445 ;
      RECT 586.14 0.155 586.4 8.665 ;
      RECT 586.65 0.155 586.91 8.665 ;
      RECT 585.63 0 585.89 11.315 ;
      RECT 586.005 74.11 586.365 74.84 ;
      RECT 586.575 74.11 586.775 74.84 ;
      RECT 587.16 0.52 587.42 9.955 ;
      RECT 587.23 74.11 587.43 74.84 ;
      RECT 587.64 74.11 588 74.84 ;
      RECT 588.295 74.11 588.495 74.84 ;
      RECT 588.79 74.11 589.15 74.84 ;
      RECT 589.2 0.3 589.46 8.7 ;
      RECT 589.36 74.11 589.56 74.84 ;
      RECT 590.015 74.11 590.215 74.84 ;
      RECT 589.71 0.18 590.48 0.88 ;
      RECT 590.425 74.11 590.785 74.84 ;
      RECT 590.995 74.11 591.195 74.84 ;
      RECT 591.65 74.11 591.85 74.84 ;
      RECT 591.905 0 592.165 6.28 ;
      RECT 592.06 74.11 592.42 74.84 ;
      RECT 592.715 74.11 592.915 74.84 ;
      RECT 593.28 0 593.54 5.57 ;
      RECT 593.21 74.11 593.57 74.84 ;
      RECT 593.78 74.11 593.98 74.84 ;
      RECT 593.79 0.3 594.05 5.235 ;
      RECT 594.3 0.52 594.56 7.78 ;
      RECT 594.435 74.11 594.635 74.84 ;
      RECT 594.845 74.11 595.205 74.84 ;
      RECT 595.15 0.52 595.41 4.315 ;
      RECT 595.415 74.11 595.615 74.84 ;
      RECT 596.07 74.11 596.27 74.84 ;
      RECT 596.325 0 596.585 2.82 ;
      RECT 596.48 74.11 596.84 74.84 ;
      RECT 597.135 74.11 597.335 74.84 ;
      RECT 597.63 74.11 597.99 74.84 ;
      RECT 598.565 0.18 599.335 0.88 ;
      RECT 598.565 0.18 598.825 12.9 ;
      RECT 599.075 0.18 599.335 12.9 ;
      RECT 597.855 0 598.115 2.82 ;
      RECT 598.2 74.11 598.4 74.84 ;
      RECT 599.585 0.155 600.355 0.445 ;
      RECT 599.585 0.155 599.845 13.21 ;
      RECT 600.095 0.155 600.355 13.21 ;
      RECT 598.855 74.11 599.055 74.84 ;
      RECT 599.265 74.11 599.625 74.84 ;
      RECT 599.835 74.11 600.035 74.84 ;
      RECT 600.49 74.11 600.69 74.84 ;
      RECT 600.9 74.11 601.26 74.84 ;
      RECT 601.555 74.11 601.755 74.84 ;
      RECT 602.05 74.11 602.41 74.84 ;
      RECT 602.29 0.52 602.55 14.115 ;
      RECT 602.62 74.11 602.82 74.84 ;
      RECT 602.8 0 603.06 13.45 ;
      RECT 603.275 74.11 603.475 74.84 ;
      RECT 603.82 0.155 604.59 0.445 ;
      RECT 603.82 0.155 604.08 8.665 ;
      RECT 604.33 0.155 604.59 8.665 ;
      RECT 603.31 0 603.57 11.315 ;
      RECT 603.685 74.11 604.045 74.84 ;
      RECT 604.255 74.11 604.455 74.84 ;
      RECT 604.84 0.52 605.1 9.955 ;
      RECT 604.91 74.11 605.11 74.84 ;
      RECT 605.32 74.11 605.68 74.84 ;
      RECT 605.975 74.11 606.175 74.84 ;
      RECT 606.47 74.11 606.83 74.84 ;
      RECT 606.88 0.3 607.14 8.7 ;
      RECT 607.04 74.11 607.24 74.84 ;
      RECT 607.695 74.11 607.895 74.84 ;
      RECT 607.39 0.18 608.16 0.88 ;
      RECT 608.105 74.11 608.465 74.84 ;
      RECT 608.675 74.11 608.875 74.84 ;
      RECT 609.33 74.11 609.53 74.84 ;
      RECT 609.585 0 609.845 6.28 ;
      RECT 609.74 74.11 610.1 74.84 ;
      RECT 610.395 74.11 610.595 74.84 ;
      RECT 610.96 0 611.22 5.57 ;
      RECT 610.89 74.11 611.25 74.84 ;
      RECT 611.46 74.11 611.66 74.84 ;
      RECT 611.47 0.3 611.73 5.235 ;
      RECT 611.98 0.52 612.24 7.78 ;
      RECT 612.115 74.11 612.315 74.84 ;
      RECT 612.525 74.11 612.885 74.84 ;
      RECT 612.83 0.52 613.09 4.315 ;
      RECT 613.095 74.11 613.295 74.84 ;
      RECT 613.75 74.11 613.95 74.84 ;
      RECT 614.005 0 614.265 2.82 ;
      RECT 614.16 74.11 614.52 74.84 ;
      RECT 614.815 74.11 615.015 74.84 ;
      RECT 615.31 74.11 615.67 74.84 ;
      RECT 616.245 0.18 617.015 0.88 ;
      RECT 616.245 0.18 616.505 12.9 ;
      RECT 616.755 0.18 617.015 12.9 ;
      RECT 615.535 0 615.795 2.82 ;
      RECT 615.88 74.11 616.08 74.84 ;
      RECT 617.265 0.155 618.035 0.445 ;
      RECT 617.265 0.155 617.525 13.21 ;
      RECT 617.775 0.155 618.035 13.21 ;
      RECT 616.535 74.11 616.735 74.84 ;
      RECT 616.945 74.11 617.305 74.84 ;
      RECT 617.515 74.11 617.715 74.84 ;
      RECT 618.17 74.11 618.37 74.84 ;
      RECT 618.58 74.11 618.94 74.84 ;
      RECT 619.235 74.11 619.435 74.84 ;
      RECT 619.73 74.11 620.09 74.84 ;
      RECT 619.97 0.52 620.23 14.115 ;
      RECT 620.3 74.11 620.5 74.84 ;
      RECT 620.48 0 620.74 13.45 ;
      RECT 620.955 74.11 621.155 74.84 ;
      RECT 621.5 0.155 622.27 0.445 ;
      RECT 621.5 0.155 621.76 8.665 ;
      RECT 622.01 0.155 622.27 8.665 ;
      RECT 620.99 0 621.25 11.315 ;
      RECT 621.365 74.11 621.725 74.84 ;
      RECT 621.935 74.11 622.135 74.84 ;
      RECT 622.52 0.52 622.78 9.955 ;
      RECT 622.59 74.11 622.79 74.84 ;
      RECT 623 74.11 623.36 74.84 ;
      RECT 623.655 74.11 623.855 74.84 ;
      RECT 624.15 74.11 624.51 74.84 ;
      RECT 624.56 0.3 624.82 8.7 ;
      RECT 624.72 74.11 624.92 74.84 ;
      RECT 625.375 74.11 625.575 74.84 ;
      RECT 625.07 0.18 625.84 0.88 ;
      RECT 625.785 74.11 626.145 74.84 ;
      RECT 626.355 74.11 626.555 74.84 ;
      RECT 627.01 74.11 627.21 74.84 ;
      RECT 627.265 0 627.525 6.28 ;
      RECT 627.42 74.11 627.78 74.84 ;
      RECT 628.075 74.11 628.275 74.84 ;
      RECT 628.64 0 628.9 5.57 ;
      RECT 628.57 74.11 628.93 74.84 ;
      RECT 629.14 74.11 629.34 74.84 ;
      RECT 629.15 0.3 629.41 5.235 ;
      RECT 629.66 0.52 629.92 7.78 ;
      RECT 629.795 74.11 629.995 74.84 ;
      RECT 630.205 74.11 630.565 74.84 ;
      RECT 630.51 0.52 630.77 4.315 ;
      RECT 630.775 74.11 630.975 74.84 ;
      RECT 631.43 74.11 631.63 74.84 ;
      RECT 631.685 0 631.945 2.82 ;
      RECT 631.84 74.11 632.2 74.84 ;
      RECT 632.495 74.11 632.695 74.84 ;
      RECT 632.99 74.11 633.35 74.84 ;
      RECT 633.925 0.18 634.695 0.88 ;
      RECT 633.925 0.18 634.185 12.9 ;
      RECT 634.435 0.18 634.695 12.9 ;
      RECT 633.215 0 633.475 2.82 ;
      RECT 633.56 74.11 633.76 74.84 ;
      RECT 634.945 0.155 635.715 0.445 ;
      RECT 634.945 0.155 635.205 13.21 ;
      RECT 635.455 0.155 635.715 13.21 ;
      RECT 634.215 74.11 634.415 74.84 ;
      RECT 634.625 74.11 634.985 74.84 ;
      RECT 635.195 74.11 635.395 74.84 ;
      RECT 635.85 74.11 636.05 74.84 ;
      RECT 636.26 74.11 636.62 74.84 ;
      RECT 636.915 74.11 637.115 74.84 ;
      RECT 637.41 74.11 637.77 74.84 ;
      RECT 637.65 0.52 637.91 14.115 ;
      RECT 637.98 74.11 638.18 74.84 ;
      RECT 638.16 0 638.42 13.45 ;
      RECT 638.635 74.11 638.835 74.84 ;
      RECT 639.18 0.155 639.95 0.445 ;
      RECT 639.18 0.155 639.44 8.665 ;
      RECT 639.69 0.155 639.95 8.665 ;
      RECT 638.67 0 638.93 11.315 ;
      RECT 639.045 74.11 639.405 74.84 ;
      RECT 639.615 74.11 639.815 74.84 ;
      RECT 640.2 0.52 640.46 9.955 ;
      RECT 640.27 74.11 640.47 74.84 ;
      RECT 640.68 74.11 641.04 74.84 ;
      RECT 641.335 74.11 641.535 74.84 ;
      RECT 641.83 74.11 642.19 74.84 ;
      RECT 642.24 0.3 642.5 8.7 ;
      RECT 642.4 74.11 642.6 74.84 ;
      RECT 643.055 74.11 643.255 74.84 ;
      RECT 642.75 0.18 643.52 0.88 ;
      RECT 643.465 74.11 643.825 74.84 ;
      RECT 644.035 74.11 644.235 74.84 ;
      RECT 644.69 74.11 644.89 74.84 ;
      RECT 644.945 0 645.205 6.28 ;
      RECT 645.1 74.11 645.46 74.84 ;
      RECT 645.755 74.11 645.955 74.84 ;
      RECT 646.32 0 646.58 5.57 ;
      RECT 646.25 74.11 646.61 74.84 ;
      RECT 646.82 74.11 647.02 74.84 ;
      RECT 646.83 0.3 647.09 5.235 ;
      RECT 647.34 0.52 647.6 7.78 ;
      RECT 647.475 74.11 647.675 74.84 ;
      RECT 647.885 74.11 648.245 74.84 ;
      RECT 648.19 0.52 648.45 4.315 ;
      RECT 648.455 74.11 648.655 74.84 ;
      RECT 649.11 74.11 649.31 74.84 ;
      RECT 649.365 0 649.625 2.82 ;
      RECT 649.52 74.11 649.88 74.84 ;
      RECT 650.175 74.11 650.375 74.84 ;
      RECT 650.67 74.11 651.03 74.84 ;
      RECT 651.605 0.18 652.375 0.88 ;
      RECT 651.605 0.18 651.865 12.9 ;
      RECT 652.115 0.18 652.375 12.9 ;
      RECT 650.895 0 651.155 2.82 ;
      RECT 651.24 74.11 651.44 74.84 ;
      RECT 652.625 0.155 653.395 0.445 ;
      RECT 652.625 0.155 652.885 13.21 ;
      RECT 653.135 0.155 653.395 13.21 ;
      RECT 651.895 74.11 652.095 74.84 ;
      RECT 652.305 74.11 652.665 74.84 ;
      RECT 652.875 74.11 653.075 74.84 ;
      RECT 653.53 74.11 653.73 74.84 ;
      RECT 653.94 74.11 654.3 74.84 ;
      RECT 654.595 74.11 654.795 74.84 ;
      RECT 655.09 74.11 655.45 74.84 ;
      RECT 655.33 0.52 655.59 14.115 ;
      RECT 655.66 74.11 655.86 74.84 ;
      RECT 655.84 0 656.1 13.45 ;
      RECT 656.315 74.11 656.515 74.84 ;
      RECT 656.86 0.155 657.63 0.445 ;
      RECT 656.86 0.155 657.12 8.665 ;
      RECT 657.37 0.155 657.63 8.665 ;
      RECT 656.35 0 656.61 11.315 ;
      RECT 656.725 74.11 657.085 74.84 ;
      RECT 657.295 74.11 657.495 74.84 ;
      RECT 657.88 0.52 658.14 9.955 ;
      RECT 657.95 74.11 658.15 74.84 ;
      RECT 658.36 74.11 658.72 74.84 ;
      RECT 659.015 74.11 659.215 74.84 ;
      RECT 659.51 74.11 659.87 74.84 ;
      RECT 659.92 0.3 660.18 8.7 ;
      RECT 660.08 74.11 660.28 74.84 ;
      RECT 660.735 74.11 660.935 74.84 ;
      RECT 660.43 0.18 661.2 0.88 ;
      RECT 661.145 74.11 661.505 74.84 ;
      RECT 661.715 74.11 661.915 74.84 ;
      RECT 662.37 74.11 662.57 74.84 ;
      RECT 662.625 0 662.885 6.28 ;
      RECT 662.78 74.11 663.14 74.84 ;
      RECT 663.435 74.11 663.635 74.84 ;
      RECT 664 0 664.26 5.57 ;
      RECT 663.93 74.11 664.29 74.84 ;
      RECT 664.5 74.11 664.7 74.84 ;
      RECT 664.51 0.3 664.77 5.235 ;
      RECT 665.02 0.52 665.28 7.78 ;
      RECT 665.155 74.11 665.355 74.84 ;
      RECT 665.565 74.11 665.925 74.84 ;
      RECT 665.87 0.52 666.13 4.315 ;
      RECT 666.135 74.11 666.335 74.84 ;
      RECT 666.79 74.11 666.99 74.84 ;
      RECT 667.045 0 667.305 2.82 ;
      RECT 667.2 74.11 667.56 74.84 ;
      RECT 667.855 74.11 668.055 74.84 ;
      RECT 668.35 74.11 668.71 74.84 ;
      RECT 669.285 0.18 670.055 0.88 ;
      RECT 669.285 0.18 669.545 12.9 ;
      RECT 669.795 0.18 670.055 12.9 ;
      RECT 668.575 0 668.835 2.82 ;
      RECT 668.92 74.11 669.12 74.84 ;
      RECT 670.305 0.155 671.075 0.445 ;
      RECT 670.305 0.155 670.565 13.21 ;
      RECT 670.815 0.155 671.075 13.21 ;
      RECT 669.575 74.11 669.775 74.84 ;
      RECT 669.985 74.11 670.345 74.84 ;
      RECT 670.555 74.11 670.755 74.84 ;
      RECT 671.21 74.11 671.41 74.84 ;
      RECT 671.62 74.11 671.98 74.84 ;
      RECT 672.275 74.11 672.475 74.84 ;
      RECT 672.77 74.11 673.13 74.84 ;
      RECT 673.01 0.52 673.27 14.115 ;
      RECT 673.34 74.11 673.54 74.84 ;
      RECT 673.52 0 673.78 13.45 ;
      RECT 673.995 74.11 674.195 74.84 ;
      RECT 674.54 0.155 675.31 0.445 ;
      RECT 674.54 0.155 674.8 8.665 ;
      RECT 675.05 0.155 675.31 8.665 ;
      RECT 674.03 0 674.29 11.315 ;
      RECT 674.405 74.11 674.765 74.84 ;
      RECT 674.975 74.11 675.175 74.84 ;
      RECT 675.56 0.52 675.82 9.955 ;
      RECT 675.63 74.11 675.83 74.84 ;
      RECT 676.04 74.11 676.4 74.84 ;
      RECT 676.695 74.11 676.895 74.84 ;
      RECT 677.19 74.11 677.55 74.84 ;
      RECT 677.6 0.3 677.86 8.7 ;
      RECT 677.76 74.11 677.96 74.84 ;
      RECT 678.415 74.11 678.615 74.84 ;
      RECT 678.11 0.18 678.88 0.88 ;
      RECT 678.825 74.11 679.185 74.84 ;
      RECT 679.395 74.11 679.595 74.84 ;
      RECT 680.05 74.11 680.25 74.84 ;
      RECT 680.305 0 680.565 6.28 ;
      RECT 680.46 74.11 680.82 74.84 ;
      RECT 681.115 74.11 681.315 74.84 ;
      RECT 681.68 0 681.94 5.57 ;
      RECT 681.61 74.11 681.97 74.84 ;
      RECT 682.18 74.11 682.38 74.84 ;
      RECT 682.19 0.3 682.45 5.235 ;
      RECT 682.7 0.52 682.96 7.78 ;
      RECT 682.835 74.11 683.035 74.84 ;
      RECT 683.245 74.11 683.605 74.84 ;
      RECT 683.55 0.52 683.81 4.315 ;
      RECT 683.815 74.11 684.015 74.84 ;
      RECT 684.47 74.11 684.67 74.84 ;
      RECT 684.725 0 684.985 2.82 ;
      RECT 684.88 74.11 685.24 74.84 ;
      RECT 685.535 74.11 685.735 74.84 ;
      RECT 686.03 74.11 686.39 74.84 ;
      RECT 686.965 0.18 687.735 0.88 ;
      RECT 686.965 0.18 687.225 12.9 ;
      RECT 687.475 0.18 687.735 12.9 ;
      RECT 686.255 0 686.515 2.82 ;
      RECT 686.6 74.11 686.8 74.84 ;
      RECT 687.985 0.155 688.755 0.445 ;
      RECT 687.985 0.155 688.245 13.21 ;
      RECT 688.495 0.155 688.755 13.21 ;
      RECT 687.255 74.11 687.455 74.84 ;
      RECT 687.665 74.11 688.025 74.84 ;
      RECT 688.235 74.11 688.435 74.84 ;
      RECT 688.89 74.11 689.09 74.84 ;
      RECT 689.3 74.11 689.66 74.84 ;
      RECT 689.955 74.11 690.155 74.84 ;
      RECT 690.45 74.11 690.81 74.84 ;
      RECT 690.69 0.52 690.95 14.115 ;
      RECT 691.02 74.11 691.22 74.84 ;
      RECT 691.2 0 691.46 13.45 ;
      RECT 691.675 74.11 691.875 74.84 ;
      RECT 692.22 0.155 692.99 0.445 ;
      RECT 692.22 0.155 692.48 8.665 ;
      RECT 692.73 0.155 692.99 8.665 ;
      RECT 691.71 0 691.97 11.315 ;
      RECT 692.085 74.11 692.445 74.84 ;
      RECT 692.655 74.11 692.855 74.84 ;
      RECT 693.24 0.52 693.5 9.955 ;
      RECT 693.31 74.11 693.51 74.84 ;
      RECT 693.72 74.11 694.08 74.84 ;
      RECT 694.375 74.11 694.575 74.84 ;
      RECT 694.87 74.11 695.23 74.84 ;
      RECT 695.28 0.3 695.54 8.7 ;
      RECT 695.44 74.11 695.64 74.84 ;
      RECT 696.095 74.11 696.295 74.84 ;
      RECT 695.79 0.18 696.56 0.88 ;
      RECT 696.505 74.11 696.865 74.84 ;
      RECT 697.075 74.11 697.275 74.84 ;
      RECT 697.73 74.11 697.93 74.84 ;
      RECT 697.985 0 698.245 6.28 ;
      RECT 698.14 74.11 698.5 74.84 ;
      RECT 698.795 74.11 698.995 74.84 ;
      RECT 699.36 0 699.62 5.57 ;
      RECT 699.29 74.11 699.65 74.84 ;
      RECT 699.86 74.11 700.06 74.84 ;
      RECT 699.87 0.3 700.13 5.235 ;
      RECT 700.38 0.52 700.64 7.78 ;
      RECT 700.515 74.11 700.715 74.84 ;
      RECT 700.925 74.11 701.285 74.84 ;
      RECT 701.495 74.11 701.695 74.84 ;
      RECT 702.32 53.41 702.52 74.84 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 426 0 427.78 74.87 ;
      RECT 443.68 0 445.46 74.87 ;
      RECT 461.36 0 463.14 74.87 ;
      RECT 479.04 0 480.82 74.87 ;
      RECT 496.72 0 498.5 74.87 ;
      RECT 514.4 0 516.18 74.87 ;
      RECT 532.08 0 533.86 74.87 ;
      RECT 549.76 0 551.54 74.87 ;
      RECT 567.44 0 569.22 74.87 ;
      RECT 585.12 0 586.9 74.87 ;
      RECT 602.8 0 604.58 74.87 ;
      RECT 620.48 0 622.26 74.87 ;
      RECT 638.16 0 639.94 74.87 ;
      RECT 655.84 0 657.62 74.87 ;
      RECT 673.52 0 675.3 74.87 ;
      RECT 691.2 0 692.98 74.87 ;
      RECT 284.74 0 315.425 74.87 ;
      RECT 327.425 0 332.765 74.87 ;
      RECT 335.585 0 335.825 74.87 ;
      RECT 356.795 0 365.715 74.87 ;
      RECT 367.005 0 367.245 74.87 ;
      RECT 370.065 0 375.405 74.87 ;
      RECT 377.195 0 386.625 74.87 ;
      RECT 428.56 0 434.92 74.87 ;
      RECT 446.24 0 452.6 74.87 ;
      RECT 463.92 0 470.28 74.87 ;
      RECT 481.6 0 487.96 74.87 ;
      RECT 499.28 0 505.64 74.87 ;
      RECT 516.96 0 523.32 74.87 ;
      RECT 534.64 0 541 74.87 ;
      RECT 552.32 0 558.68 74.87 ;
      RECT 570 0 576.36 74.87 ;
      RECT 587.68 0 594.04 74.87 ;
      RECT 605.36 0 611.72 74.87 ;
      RECT 623.04 0 629.4 74.87 ;
      RECT 640.72 0 647.08 74.87 ;
      RECT 658.4 0 664.76 74.87 ;
      RECT 676.08 0 682.44 74.87 ;
      RECT 693.76 0 700.12 74.87 ;
      RECT 0 0 1.93 74.87 ;
      RECT 2.71 0 9.07 74.87 ;
      RECT 2.7 0.3 9.07 74.87 ;
      RECT 9.85 0 11.63 74.87 ;
      RECT 9.84 0.155 11.63 74.87 ;
      RECT 12.4 0 18.76 74.87 ;
      RECT 20.39 0 26.75 74.87 ;
      RECT 20.38 0.3 26.75 74.87 ;
      RECT 27.53 0 29.31 74.87 ;
      RECT 27.52 0.155 29.31 74.87 ;
      RECT 30.08 0 36.44 74.87 ;
      RECT 38.07 0 44.43 74.87 ;
      RECT 38.06 0.3 44.43 74.87 ;
      RECT 45.21 0 46.99 74.87 ;
      RECT 45.2 0.155 46.99 74.87 ;
      RECT 47.76 0 54.12 74.87 ;
      RECT 55.75 0 62.11 74.87 ;
      RECT 55.74 0.3 62.11 74.87 ;
      RECT 62.89 0 64.67 74.87 ;
      RECT 62.88 0.155 64.67 74.87 ;
      RECT 65.44 0 71.8 74.87 ;
      RECT 73.43 0 79.79 74.87 ;
      RECT 73.42 0.3 79.79 74.87 ;
      RECT 80.57 0 82.35 74.87 ;
      RECT 80.56 0.155 82.35 74.87 ;
      RECT 83.12 0 89.48 74.87 ;
      RECT 91.11 0 97.47 74.87 ;
      RECT 91.1 0.3 97.47 74.87 ;
      RECT 98.25 0 100.03 74.87 ;
      RECT 98.24 0.155 100.03 74.87 ;
      RECT 100.8 0 107.16 74.87 ;
      RECT 108.79 0 115.15 74.87 ;
      RECT 108.78 0.3 115.15 74.87 ;
      RECT 115.93 0 117.71 74.87 ;
      RECT 115.92 0.155 117.71 74.87 ;
      RECT 118.48 0 124.84 74.87 ;
      RECT 126.47 0 132.83 74.87 ;
      RECT 126.46 0.3 132.83 74.87 ;
      RECT 133.61 0 135.39 74.87 ;
      RECT 133.6 0.155 135.39 74.87 ;
      RECT 136.16 0 142.52 74.87 ;
      RECT 144.15 0 150.51 74.87 ;
      RECT 144.14 0.3 150.51 74.87 ;
      RECT 151.29 0 153.07 74.87 ;
      RECT 151.28 0.155 153.07 74.87 ;
      RECT 153.84 0 160.2 74.87 ;
      RECT 161.83 0 168.19 74.87 ;
      RECT 161.82 0.3 168.19 74.87 ;
      RECT 168.97 0 170.75 74.87 ;
      RECT 168.96 0.155 170.75 74.87 ;
      RECT 171.52 0 177.88 74.87 ;
      RECT 179.51 0 185.87 74.87 ;
      RECT 179.5 0.3 185.87 74.87 ;
      RECT 186.65 0 188.43 74.87 ;
      RECT 186.64 0.155 188.43 74.87 ;
      RECT 189.2 0 195.56 74.87 ;
      RECT 197.19 0 203.55 74.87 ;
      RECT 197.18 0.3 203.55 74.87 ;
      RECT 204.33 0 206.11 74.87 ;
      RECT 204.32 0.155 206.11 74.87 ;
      RECT 206.88 0 213.24 74.87 ;
      RECT 214.87 0 221.23 74.87 ;
      RECT 214.86 0.3 221.23 74.87 ;
      RECT 222.01 0 223.79 74.87 ;
      RECT 222 0.155 223.79 74.87 ;
      RECT 224.56 0 230.92 74.87 ;
      RECT 232.55 0 238.91 74.87 ;
      RECT 232.54 0.3 238.91 74.87 ;
      RECT 239.69 0 241.47 74.87 ;
      RECT 239.68 0.155 241.47 74.87 ;
      RECT 242.24 0 248.6 74.87 ;
      RECT 250.23 0 256.59 74.87 ;
      RECT 250.22 0.3 256.59 74.87 ;
      RECT 257.37 0 259.15 74.87 ;
      RECT 257.36 0.155 259.15 74.87 ;
      RECT 259.92 0 266.28 74.87 ;
      RECT 267.91 0 274.27 74.87 ;
      RECT 267.9 0.3 274.27 74.87 ;
      RECT 275.05 0 276.83 74.87 ;
      RECT 275.04 0.155 276.83 74.87 ;
      RECT 277.6 0 283.96 74.87 ;
      RECT 284.74 0.18 315.435 74.87 ;
      RECT 316.205 0 325.635 74.87 ;
      RECT 316.195 0.3 325.635 74.87 ;
      RECT 326.395 0 326.655 74.87 ;
      RECT 327.415 0.3 332.775 74.87 ;
      RECT 334.045 0 334.305 74.87 ;
      RECT 335.575 0.3 335.835 74.87 ;
      RECT 337.115 0 346.035 74.87 ;
      RECT 337.105 0.3 346.035 74.87 ;
      RECT 346.795 0 347.055 74.87 ;
      RECT 347.815 0 355.015 74.87 ;
      RECT 355.775 0 356.035 74.87 ;
      RECT 356.795 0.3 365.725 74.87 ;
      RECT 366.995 0.3 367.255 74.87 ;
      RECT 368.525 0 368.785 74.87 ;
      RECT 370.055 0.3 375.415 74.87 ;
      RECT 376.175 0 376.435 74.87 ;
      RECT 377.195 0.3 386.635 74.87 ;
      RECT 387.405 0 418.09 74.87 ;
      RECT 387.395 0.18 418.09 74.87 ;
      RECT 418.87 0 425.23 74.87 ;
      RECT 426 0.155 427.79 74.87 ;
      RECT 428.56 0.3 434.93 74.87 ;
      RECT 436.55 0 442.91 74.87 ;
      RECT 443.68 0.155 445.47 74.87 ;
      RECT 446.24 0.3 452.61 74.87 ;
      RECT 454.23 0 460.59 74.87 ;
      RECT 461.36 0.155 463.15 74.87 ;
      RECT 463.92 0.3 470.29 74.87 ;
      RECT 471.91 0 478.27 74.87 ;
      RECT 479.04 0.155 480.83 74.87 ;
      RECT 481.6 0.3 487.97 74.87 ;
      RECT 489.59 0 495.95 74.87 ;
      RECT 496.72 0.155 498.51 74.87 ;
      RECT 499.28 0.3 505.65 74.87 ;
      RECT 507.27 0 513.63 74.87 ;
      RECT 514.4 0.155 516.19 74.87 ;
      RECT 516.96 0.3 523.33 74.87 ;
      RECT 524.95 0 531.31 74.87 ;
      RECT 532.08 0.155 533.87 74.87 ;
      RECT 534.64 0.3 541.01 74.87 ;
      RECT 542.63 0 548.99 74.87 ;
      RECT 549.76 0.155 551.55 74.87 ;
      RECT 552.32 0.3 558.69 74.87 ;
      RECT 560.31 0 566.67 74.87 ;
      RECT 567.44 0.155 569.23 74.87 ;
      RECT 570 0.3 576.37 74.87 ;
      RECT 577.99 0 584.35 74.87 ;
      RECT 585.12 0.155 586.91 74.87 ;
      RECT 587.68 0.3 594.05 74.87 ;
      RECT 595.67 0 602.03 74.87 ;
      RECT 602.8 0.155 604.59 74.87 ;
      RECT 605.36 0.3 611.73 74.87 ;
      RECT 613.35 0 619.71 74.87 ;
      RECT 620.48 0.155 622.27 74.87 ;
      RECT 623.04 0.3 629.41 74.87 ;
      RECT 631.03 0 637.39 74.87 ;
      RECT 638.16 0.155 639.95 74.87 ;
      RECT 640.72 0.3 647.09 74.87 ;
      RECT 648.71 0 655.07 74.87 ;
      RECT 655.84 0.155 657.63 74.87 ;
      RECT 658.4 0.3 664.77 74.87 ;
      RECT 666.39 0 672.75 74.87 ;
      RECT 673.52 0.155 675.31 74.87 ;
      RECT 676.08 0.3 682.45 74.87 ;
      RECT 684.07 0 690.43 74.87 ;
      RECT 691.2 0.155 692.99 74.87 ;
      RECT 693.76 0.3 700.13 74.87 ;
      RECT 700.9 0 702.83 74.87 ;
      RECT 0 0.52 702.83 74.87 ;
    LAYER Metal3 ;
      RECT 0 0 702.83 74.87 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 0 47.305 14.725 53.15 ;
      RECT 0 0 5.885 74.87 ;
      RECT 10.825 0 14.725 74.87 ;
      RECT 19.665 47.305 32.405 53.15 ;
      RECT 19.665 0 23.565 74.87 ;
      RECT 28.505 0 32.405 74.87 ;
      RECT 37.345 47.305 50.085 53.15 ;
      RECT 37.345 0 41.245 74.87 ;
      RECT 46.185 0 50.085 74.87 ;
      RECT 55.025 47.305 67.765 53.15 ;
      RECT 55.025 0 58.925 74.87 ;
      RECT 63.865 0 67.765 74.87 ;
      RECT 72.705 47.305 85.445 53.15 ;
      RECT 72.705 0 76.605 74.87 ;
      RECT 81.545 0 85.445 74.87 ;
      RECT 90.385 47.305 103.125 53.15 ;
      RECT 90.385 0 94.285 74.87 ;
      RECT 99.225 0 103.125 74.87 ;
      RECT 108.065 47.305 120.805 53.15 ;
      RECT 108.065 0 111.965 74.87 ;
      RECT 116.905 0 120.805 74.87 ;
      RECT 125.745 47.305 138.485 53.15 ;
      RECT 125.745 0 129.645 74.87 ;
      RECT 134.585 0 138.485 74.87 ;
      RECT 143.425 47.305 156.165 53.15 ;
      RECT 143.425 0 147.325 74.87 ;
      RECT 152.265 0 156.165 74.87 ;
      RECT 161.105 47.305 173.845 53.15 ;
      RECT 161.105 0 165.005 74.87 ;
      RECT 169.945 0 173.845 74.87 ;
      RECT 178.785 47.305 191.525 53.15 ;
      RECT 178.785 0 182.685 74.87 ;
      RECT 187.625 0 191.525 74.87 ;
      RECT 196.465 47.305 209.205 53.15 ;
      RECT 196.465 0 200.365 74.87 ;
      RECT 205.305 0 209.205 74.87 ;
      RECT 214.145 47.305 226.885 53.15 ;
      RECT 214.145 0 218.045 74.87 ;
      RECT 222.985 0 226.885 74.87 ;
      RECT 231.825 47.305 244.565 53.15 ;
      RECT 231.825 0 235.725 74.87 ;
      RECT 240.665 0 244.565 74.87 ;
      RECT 249.505 47.305 262.245 53.15 ;
      RECT 249.505 0 253.405 74.87 ;
      RECT 258.345 0 262.245 74.87 ;
      RECT 267.185 47.305 279.925 53.15 ;
      RECT 267.185 0 271.085 74.87 ;
      RECT 276.025 0 279.925 74.87 ;
      RECT 284.865 0 311.125 74.87 ;
      RECT 314.455 0 316.275 74.87 ;
      RECT 319.605 0 321.425 74.87 ;
      RECT 324.755 0 326.575 74.87 ;
      RECT 329.905 0 331.725 74.87 ;
      RECT 335.055 0 336.875 74.87 ;
      RECT 340.205 0 342.025 74.87 ;
      RECT 345.355 0 347.175 74.87 ;
      RECT 350.505 0 352.325 74.87 ;
      RECT 355.655 0 357.475 74.87 ;
      RECT 360.805 0 362.625 74.87 ;
      RECT 365.955 0 367.775 74.87 ;
      RECT 371.105 0 372.925 74.87 ;
      RECT 376.255 0 378.075 74.87 ;
      RECT 422.905 47.305 435.645 53.15 ;
      RECT 422.905 0 426.805 74.87 ;
      RECT 431.745 0 435.645 74.87 ;
      RECT 440.585 47.305 453.325 53.15 ;
      RECT 440.585 0 444.485 74.87 ;
      RECT 449.425 0 453.325 74.87 ;
      RECT 458.265 47.305 471.005 53.15 ;
      RECT 458.265 0 462.165 74.87 ;
      RECT 467.105 0 471.005 74.87 ;
      RECT 475.945 47.305 488.685 53.15 ;
      RECT 475.945 0 479.845 74.87 ;
      RECT 484.785 0 488.685 74.87 ;
      RECT 493.625 47.305 506.365 53.15 ;
      RECT 493.625 0 497.525 74.87 ;
      RECT 502.465 0 506.365 74.87 ;
      RECT 511.305 47.305 524.045 53.15 ;
      RECT 511.305 0 515.205 74.87 ;
      RECT 520.145 0 524.045 74.87 ;
      RECT 528.985 47.305 541.725 53.15 ;
      RECT 528.985 0 532.885 74.87 ;
      RECT 537.825 0 541.725 74.87 ;
      RECT 546.665 47.305 559.405 53.15 ;
      RECT 546.665 0 550.565 74.87 ;
      RECT 555.505 0 559.405 74.87 ;
      RECT 564.345 47.305 577.085 53.15 ;
      RECT 564.345 0 568.245 74.87 ;
      RECT 573.185 0 577.085 74.87 ;
      RECT 582.025 47.305 594.765 53.15 ;
      RECT 582.025 0 585.925 74.87 ;
      RECT 590.865 0 594.765 74.87 ;
      RECT 599.705 47.305 612.445 53.15 ;
      RECT 599.705 0 603.605 74.87 ;
      RECT 608.545 0 612.445 74.87 ;
      RECT 617.385 47.305 630.125 53.15 ;
      RECT 617.385 0 621.285 74.87 ;
      RECT 626.225 0 630.125 74.87 ;
      RECT 635.065 47.305 647.805 53.15 ;
      RECT 635.065 0 638.965 74.87 ;
      RECT 643.905 0 647.805 74.87 ;
      RECT 652.745 47.305 665.485 53.15 ;
      RECT 652.745 0 656.645 74.87 ;
      RECT 661.585 0 665.485 74.87 ;
      RECT 670.425 47.305 683.165 53.15 ;
      RECT 670.425 0 674.325 74.87 ;
      RECT 679.265 0 683.165 74.87 ;
      RECT 688.105 47.305 702.83 53.15 ;
      RECT 688.105 0 692.005 74.87 ;
      RECT 696.945 0 702.83 74.87 ;
      RECT 381.405 0 383.225 74.87 ;
      RECT 386.555 0 388.375 74.87 ;
      RECT 391.705 0 417.965 74.87 ;
  END
END RM_IHPSG13_2P_64x32_c2

END LIBRARY
