************************************************************************
* 
* Copyright 2023 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
************************************************************************
* auCdl Netlist:
* 
* Library Name:  sg13g2_stdcell
* Top Cell Name: sg13g2_stdcell_allcells
* View Name:     schematic
* Netlisted on:  Mar 29 14:17:55 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and2_1 A B VSS VDD X
*.PININFO A:B B:B VDD:B VSS:B X:B
MX0 a_56_136_ A a_143_136_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 VSS a_56_136_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 a_143_136_ B VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 a_56_136_ B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 VDD a_56_136_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 VDD A a_56_136_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and3_1 A B C VSS VDD X
*.PININFO A:B B:B C:B VDD:B VSS:B X:B
MX0 a_233_136_ C VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 VSS a_27_398_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_27_398_ A a_121_136_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX6 a_121_136_ B a_233_136_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 VDD B a_27_398_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 VDD a_27_398_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX4 a_27_398_ A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 a_27_398_ C VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and4_1 A B C D VSS VDD X
*.PININFO A:B B:B C:B D:B VDD:B VSS:B X:B
MX0 a_96_74_ A a_179_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 a_257_74_ C a_335_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX4 VSS a_96_74_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 a_335_74_ D VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 a_179_74_ B a_257_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 VDD a_96_74_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 VDD A a_96_74_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 VDD C a_96_74_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX6 a_96_74_ B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX9 a_96_74_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_1 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_16
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_16 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=4.44u l=130.00n ng=6
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=11.84u l=130.00n ng=16
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=17.92u l=130.00n ng=16
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=6.72u l=130.00n ng=6
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_2 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=1.48u l=130.00n ng=2
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=2.24u l=130.00n ng=2
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_4 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=2.96u l=130.00n ng=4
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=4.48u l=130.00n ng=4
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=1.68u l=130.00n ng=2
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_8 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=2.22u l=130.00n ng=3
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=5.92u l=130.00n ng=8
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=8.96u l=130.00n ng=8
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=3.36u l=130.00n ng=3
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dfrbp_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dfrbp_2 CLK D RESET_B VSS VDD Q Q_N
*.PININFO CLK:B D:B Q:B Q_N:B RESET_B:B VDD:B VSS:B
MX28 VDD D a_70_74_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX15 a_1755_389_ a_1800_291_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX20 a_1586_149_ a_818_418_ a_1755_389_ VDD sg13_lv_pmos m=1 w=420.00n 
+ l=130.00n ng=1
MX19 VDD a_331_392_ a_683_485_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX37 a_683_485_ a_728_331_ a_298_294_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX23 VDD CLK a_728_331_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 a_1800_291_ a_1586_149_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX35 VDD RESET_B a_1800_291_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX5 a_818_418_ a_728_331_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX22 a_298_294_ a_818_418_ a_70_74_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX33 a_331_392_ a_728_331_ a_1586_149_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX32 VDD a_298_294_ a_331_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 a_298_294_ RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX27 a_70_74_ RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX31 Q_N a_1586_149_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX13 VDD a_1586_149_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX24 VDD a_1586_149_ a_2363_352_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX25 Q a_2363_352_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 VDD a_2363_352_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX30 VSS RESET_B a_536_81_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX34 a_536_81_ a_331_392_ a_614_81_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX29 a_298_294_ a_818_418_ a_614_81_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX0 a_156_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX17 a_70_74_ D a_156_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX36 a_1499_149_ a_728_331_ a_1586_149_ VSS sg13_lv_nmos m=1 w=420.00n 
+ l=130.00n ng=1
MX11 a_1499_149_ a_1800_291_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX21 a_1974_74_ a_1586_149_ a_1800_291_ VSS sg13_lv_nmos m=1 w=420.00n 
+ l=130.00n ng=1
MX14 VSS RESET_B a_1974_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX12 VSS CLK a_728_331_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 a_818_418_ a_728_331_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX26 VSS a_298_294_ a_331_392_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 a_1586_149_ a_818_418_ a_331_392_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
MX1 a_70_74_ a_728_331_ a_298_294_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX18 Q_N a_1586_149_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 VSS a_1586_149_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX9 VSS a_1586_149_ a_2363_352_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX10 Q a_2363_352_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 VSS a_2363_352_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlygate4sd1_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlygate4sd1_1 A VSS VDD X
*.PININFO A:B VDD:B VSS:B X:B
MX0 VDD a_405_138_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 VDD a_28_74_ a_286_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 a_405_138_ a_286_392_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX5 a_28_74_ A VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX2 a_28_74_ A VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX3 VSS a_405_138_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 a_405_138_ a_286_392_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX7 VSS a_28_74_ a_286_392_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlygate4sd2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlygate4sd2_1 A VSS VDD X
*.PININFO A:B VDD:B VSS:B X:B
MX0 VDD a_405_138_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 VDD a_28_74_ a_288_74_ VDD sg13_lv_pmos m=1 w=1.000u l=250.00n ng=1
MX2 a_405_138_ a_288_74_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=250.00n ng=1
MX6 a_28_74_ A VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX3 VSS a_28_74_ a_288_74_ VSS sg13_lv_nmos m=1 w=420.00n l=180.00n ng=1
MX4 a_28_74_ A VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX5 VSS a_405_138_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 a_405_138_ a_288_74_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=180.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlygate4sd3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlygate4sd3_1 A VSS VDD X
*.PININFO A:B VDD:B VSS:B X:B
MX0 a_405_138_ a_289_74_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=500.0n ng=1
MX1 VDD a_405_138_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 a_28_74_ A VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX7 VDD a_28_74_ a_289_74_ VDD sg13_lv_pmos m=1 w=1.000u l=500.0n ng=1
MX2 VSS a_28_74_ a_289_74_ VSS sg13_lv_nmos m=1 w=420.00n l=500.0n ng=1
MX3 a_405_138_ a_289_74_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=500.0n ng=1
MX4 a_28_74_ A VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX5 VSS a_405_138_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_1 A VDD VSS Y
*.PININFO A:B VDD:B VSS:B Y:B
MX1 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX0 VDD A Y VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_16
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_16 A VSS VDD Y
*.PININFO A:B VDD:B VSS:B Y:B
MX30 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX29 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX27 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX21 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX19 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX9 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX31 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX28 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX26 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX25 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX24 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX23 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX20 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX15 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX14 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX13 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX4 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX0 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_2 A VDD VSS Y
*.PININFO A:B VDD:B VSS:B Y:B
MX0 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_4 A VSS VDD Y
*.PININFO A:B VDD:B VSS:B Y:B
MX0 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_8 A VSS VDD Y
*.PININFO A:B VDD:B VSS:B Y:B
MX0 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX13 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX14 VDD A Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX15 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_mux2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_mux2_1 A0 A1 S VSS VDD X
*.PININFO A0:B A1:B S:B VDD:B VSS:B X:B
MX0 a_223_368_ A0 a_304_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX2 VDD S a_223_368_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX6 a_27_112_ S VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 a_524_368_ a_27_112_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX9 VDD a_304_74_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 a_304_74_ A1 a_524_368_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX1 VSS S a_226_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 a_443_74_ a_27_112_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 VSS a_304_74_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_304_74_ A0 a_443_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 a_226_74_ A1 a_304_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 a_27_112_ S VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a21o_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a21o_1 A1 A2 B1 VSS VDD X
*.PININFO A1:B A2:B B1:B VDD:B VSS:B X:B
MX0 a_452_136_ A2 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 VSS B1 a_81_264_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX4 a_81_264_ A1 a_452_136_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX7 X a_81_264_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 a_81_264_ B1 a_364_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX3 X a_81_264_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 a_364_392_ A1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX6 VDD A2 a_364_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_mux4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_mux4_1 A0 A1 A2 A3 S0 S1 VSS VDD X
*.PININFO A0:B A1:B A2:B A3:B S0:B S1:B VDD:B VSS:B X:B
MX2 VDD A0 a_255_341_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX21 a_255_341_ S0 a_342_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX14 a_537_341_ A1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX6 a_342_74_ a_27_74_ a_537_341_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX24 VDD A2 a_763_341_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX17 a_763_341_ S0 a_846_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX20 a_1065_387_ A3 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX25 a_846_74_ a_27_74_ a_1065_387_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX16 VDD a_1338_125_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX10 a_27_74_ S0 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX11 a_1338_125_ a_1396_99_ a_846_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX5 a_342_74_ S1 a_1338_125_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX0 a_1396_99_ S1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX1 a_264_74_ a_27_74_ a_342_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 VSS A0 a_264_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX3 a_342_74_ S0 a_450_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX22 a_450_74_ A1 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX4 a_768_74_ a_27_74_ a_846_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX12 VSS A2 a_768_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX9 a_846_74_ S0 a_979_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX15 a_979_74_ A3 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX13 VSS a_1338_125_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX19 a_27_74_ S0 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX7 a_846_74_ S1 a_1338_125_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX18 a_1338_125_ a_1396_99_ a_342_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n 
+ ng=1
MX23 a_1396_99_ S1 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand2_1 A B VSS VDD Y
*.PININFO A:B B:B VDD:B VSS:B Y:B
MX0 VDD B Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_117_74_ A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS B a_117_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand2b_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand2b_1 A_N B VSS VDD Y
*.PININFO A_N:B B:B VDD:B VSS:B Y:B
MX0 Y a_27_112_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 a_27_112_ A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 VDD B Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_269_74_ a_27_112_ Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_27_112_ A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX5 VSS B a_269_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand3b_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand3b_1 A_N B C VSS VDD Y
*.PININFO A_N:B B:B C:B VDD:B VSS:B Y:B
MX0 a_27_116_ A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 VDD a_27_116_ Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 VDD C Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 a_269_78_ B a_347_78_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_347_78_ a_27_116_ Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_27_116_ A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 VSS C a_269_78_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor2_1 A B VSS VDD Y
*.PININFO A:B B:B VDD:B VSS:B Y:B
MX0 Y B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 VDD A a_116_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_116_368_ B Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor3_1 A B C VSS VDD Y
*.PININFO A:B B:B C:B VDD:B VSS:B Y:B
MX0 a_114_368_ B a_198_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 VDD A a_114_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 a_198_368_ C Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 VSS C Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor4_1 A B C D VSS VDD Y
*.PININFO A:B B:B C:B D:B VDD:B VSS:B Y:B
MX0 VDD A a_144_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 a_144_368_ B a_228_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 a_228_368_ C a_342_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 a_342_368_ D Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 VSS C Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 VSS A Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 Y D VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 Y B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or2_1 A B VDD VSS X
*.PININFO A:B B:B VDD:B VSS:B X:B
MP0 net2 B net3 VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP1 net3 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 X net2 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MN0 net2 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN1 net2 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 X net2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or3_1 A B C VSS VDD X
*.PININFO A:B B:B C:B VDD:B VSS:B X:B
MX0 a_27_74_ A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 VSS a_27_74_ X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 a_27_74_ C VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 VSS B a_27_74_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX2 VDD a_27_74_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 a_27_74_ C a_116_368_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 a_116_368_ B a_200_368_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX5 a_200_368_ A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or4_1 A B C D VDD VSS X
*.PININFO A:I B:I C:I D:I X:O VDD:B VSS:B
MN4 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN3 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 net1 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN1 net1 C VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN0 net1 D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MP4 net4 D VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP3 net3 C net4 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP2 net2 B net3 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net1 A net2 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP0 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_xnor2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_xnor2_1 A B VSS VDD Y
*.PININFO A:B B:B VDD:B VSS:B Y:B
MX0 a_376_368_ B Y VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y a_138_385_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_138_385_ B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 VDD A a_138_385_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX9 VDD A a_376_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX4 VSS B a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_112_119_ B a_138_385_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX6 VSS A a_112_119_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX7 a_293_74_ A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 a_293_74_ a_138_385_ Y VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_xor2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_xor2_1 A B VSS VDD X
*.PININFO A:B B:B VDD:B VSS:B X:B
MX0 VSS A a_194_125_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX4 a_455_87_ B X VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 X a_194_125_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 VSS A a_455_87_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX9 a_194_125_ B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 VDD A a_158_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX2 a_158_392_ B a_194_125_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX3 a_355_368_ A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 VDD B a_355_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 a_355_368_ a_194_125_ X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dfrbp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dfrbp_1 CLK D Q Q_N RESET_B VDD VSS
*.PININFO CLK:B D:B Q:B Q_N:B RESET_B:B VDD:B VSS:B
MX32 VDD D a_38_78_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX20 a_705_463_ a_319_392_ a_796_463_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX4 a_796_463_ a_841_401_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX19 a_319_392_ CLK VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX22 a_1224_74_ a_500_392_ a_1465_471_ VDD sg13_lv_pmos m=1 w=420.00n 
+ l=130.00n ng=1
MX15 a_1465_471_ a_1482_48_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX23 VDD a_1224_74_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX29 VDD a_2026_424_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 VDD a_705_463_ a_841_401_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX21 VDD RESET_B a_705_463_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX1 a_38_78_ a_500_392_ a_705_463_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX6 a_38_78_ RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX13 VDD a_319_392_ a_500_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX0 VDD RESET_B a_1482_48_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX8 a_841_401_ a_319_392_ a_1224_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX16 a_1482_48_ a_1224_74_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX26 a_2026_424_ a_1224_74_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX2 a_705_463_ a_500_392_ a_832_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX30 a_832_119_ a_841_401_ a_910_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX17 a_910_119_ RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX7 a_125_78_ RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 a_38_78_ D a_125_78_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX14 a_319_392_ CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX25 VSS RESET_B a_1624_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX9 a_1624_74_ a_1224_74_ a_1482_48_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX24 a_1224_74_ a_319_392_ a_1434_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX28 a_1434_74_ a_1482_48_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX12 VSS a_1224_74_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 VSS a_2026_424_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS a_705_463_ a_841_401_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX31 a_38_78_ a_319_392_ a_705_463_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX27 VSS a_319_392_ a_500_392_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX33 a_841_401_ a_500_392_ a_1224_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n 
+ ng=1
MX18 a_2026_424_ a_1224_74_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_sdfbbp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_sdfbbp_1 CLK D Q Q_N RESET_B SCD SCE SET_B VDD VSS
*.PININFO CLK:B D:B Q:B Q_N:B RESET_B:B SCD:B SCE:B SET_B:B VDD:B VSS:B
MX46 a_1625_93_ RESET_B VDD VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX45 a_2037_442_ a_1878_420_ a_2384_392_ VDD sg13_lv_pmos m=1 w=1.000u 
+ l=130.00n ng=1
MX44 VDD SET_B a_2037_442_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX41 VDD a_622_98_ a_877_98_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX39 VDD SCE a_341_93_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX38 a_218_464_ D a_197_119_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX33 a_1092_96_ a_622_98_ a_1221_419_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX28 a_1221_419_ a_1250_231_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX27 VDD SCE a_218_464_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX26 VDD a_2037_442_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX24 VDD a_1250_231_ a_1766_379_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX19 a_2384_392_ a_1625_93_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX17 VDD SET_B a_1250_231_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX16 a_27_464_ SCD VDD VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX15 a_622_98_ CLK VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX14 a_1250_231_ a_1092_96_ a_1580_379_ VDD sg13_lv_pmos m=1 w=840.00n 
+ l=130.00n ng=1
MX11 a_197_119_ a_877_98_ a_1092_96_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n 
+ ng=1
MX9 a_197_119_ a_341_93_ a_27_464_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n 
+ ng=1
MX8 a_2881_74_ a_2037_442_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 a_1580_379_ a_1625_93_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX6 a_1986_504_ a_2037_442_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX5 a_1878_420_ a_877_98_ a_1986_504_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX4 a_1766_379_ a_622_98_ a_1878_420_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n 
+ ng=1
MX3 VDD a_2881_74_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX47 a_2271_74_ a_1878_420_ a_2037_442_ VSS sg13_lv_nmos m=1 w=740.00n 
+ l=130.00n ng=1
MX43 a_197_119_ a_622_98_ a_1092_96_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX42 a_299_119_ a_341_93_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX40 VSS a_622_98_ a_877_98_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX37 a_1625_93_ RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX36 a_2061_74_ a_2037_442_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX35 a_1418_125_ a_1092_96_ a_1250_231_ VSS sg13_lv_nmos m=1 w=550.00n 
+ l=130.00n ng=1
MX34 VSS SCE a_341_93_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX32 VSS SET_B a_1418_125_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX31 a_1192_96_ a_1250_231_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX30 a_119_119_ SCE a_197_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX29 VSS SET_B a_2271_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX25 a_1092_96_ a_877_98_ a_1192_96_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX23 a_197_119_ D a_299_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX22 a_2881_74_ a_2037_442_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX21 a_1878_420_ a_622_98_ a_2061_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX20 VSS a_2881_74_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 VSS a_1250_231_ a_1880_119_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX13 a_622_98_ CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 VSS SCD a_119_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 a_1880_119_ a_877_98_ a_1878_420_ VSS sg13_lv_nmos m=1 w=550.00n 
+ l=130.00n ng=1
MX2 a_1250_231_ a_1625_93_ a_1418_125_ VSS sg13_lv_nmos m=1 w=550.00n 
+ l=130.00n ng=1
MX1 VSS a_2037_442_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX0 a_2037_442_ a_1625_93_ a_2271_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_lgcp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_lgcp_1 CLK GATE GCLK VDD VSS
*.PININFO CLK:B GATE:B GCLK:B VDD:B VSS:B
MX15 VDD a_315_54_ a_309_338_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX14 a_258_392_ a_309_338_ a_83_260_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX12 a_27_74_ a_83_260_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 VDD GATE a_258_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX9 a_987_393_ a_27_74_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 VDD a_987_393_ GCLK VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 a_83_260_ a_315_54_ a_484_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX4 a_315_54_ CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 VDD CLK a_987_393_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX2 a_484_508_ a_27_74_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX19 VSS a_987_393_ GCLK VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 a_984_125_ a_27_74_ a_987_393_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n 
+ ng=1
MX17 a_27_74_ a_83_260_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 VSS a_315_54_ a_309_338_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX13 a_477_124_ a_27_74_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 VSS GATE a_267_80_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 a_83_260_ a_309_338_ a_477_124_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX6 a_315_54_ CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 VSS CLK a_984_125_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX0 a_267_80_ a_315_54_ a_83_260_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_slgcp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_slgcp_1 CLK GATE GCLK SCE VDD VSS
*.PININFO CLK:B GATE:B GCLK:B SCE:B VDD:B VSS:B
MX19 GCLK a_1238_94_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX18 a_114_112_ CLKbb a_566_74_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX16 CLKbb CLKb VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX14 a_1238_94_ a_709_54_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX13 a_116_424_ SCE VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX11 a_566_74_ CLKb a_722_492_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX9 a_709_54_ a_566_74_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 CLKb CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 a_1238_94_ CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 a_722_492_ a_709_54_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX2 a_114_112_ GATE a_116_424_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX21 a_709_54_ a_566_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX20 net2 CLK VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX17 a_114_112_ SCE VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX15 a_566_74_ CLKb a_114_112_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX12 a_667_80_ a_709_54_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 a_1238_94_ a_709_54_ net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 GCLK a_1238_94_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 CLKbb CLKb VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_114_112_ GATE VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 CLKb CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX0 a_566_74_ CLKbb a_667_80_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlhq_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlhq_1 D GATE Q VDD VSS
*.PININFO D:B GATE:B Q:B VDD:B VSS:B
MX17 VDD a_386_326_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX16 a_592_149_ a_685_59_ a_419_392_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX14 a_386_326_ a_592_149_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX12 VDD D a_116_424_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX9 a_562_123_ GATE VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 VDD a_562_123_ a_685_59_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 VDD a_386_326_ a_419_392_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX3 a_229_392_ a_562_123_ a_592_149_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX1 a_229_392_ a_116_424_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX15 a_562_123_ GATE VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX13 VSS a_562_123_ a_685_59_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 a_514_149_ a_562_123_ a_592_149_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX10 VSS a_386_326_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 a_239_85_ a_116_424_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 VSS a_386_326_ a_514_149_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX5 a_386_326_ a_592_149_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 a_592_149_ a_685_59_ a_239_85_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
MX0 VSS D a_116_424_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlhr_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlhr_1 D GATE Q Q_N RESET_B VDD VSS
*.PININFO D:B GATE:B Q:B Q_N:B RESET_B:B VDD:B VSS:B
MX0 a_823_98_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 VDD a_823_98_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX15 a_642_392_ a_353_98_ a_753_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX6 a_753_508_ a_823_98_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX10 a_564_392_ a_226_104_ a_642_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX18 VDD a_27_142_ a_564_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX13 a_27_142_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 VDD GATE a_226_104_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 VDD a_1342_74_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 VDD a_642_392_ a_823_98_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX20 a_353_98_ a_226_104_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX2 a_1342_74_ a_823_98_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX12 a_823_98_ a_642_392_ a_1051_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
MX21 a_1051_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 a_642_392_ a_226_104_ a_775_124_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX14 a_775_124_ a_823_98_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX7 VSS a_823_98_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 a_571_80_ a_353_98_ a_642_392_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n 
+ ng=1
MX23 VSS a_27_142_ a_571_80_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX4 a_27_142_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX19 VSS GATE a_226_104_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 VSS a_1342_74_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 a_353_98_ a_226_104_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 a_1342_74_ a_823_98_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlhrq_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlhrq_1 D GATE Q RESET_B VDD VSS
*.PININFO D:B GATE:B Q:B RESET_B:B VDD:B VSS:B
MX19 a_769_74_ a_817_48_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX14 a_565_74_ a_363_74_ a_643_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n 
+ ng=1
MX11 VSS a_817_48_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 a_27_424_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX8 a_1045_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 a_817_48_ a_643_74_ a_1045_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
MX6 a_643_74_ a_216_424_ a_769_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX4 VSS GATE a_216_424_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS a_27_424_ a_565_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 a_363_74_ a_216_424_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 VDD a_643_74_ a_817_48_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX17 VDD a_27_424_ a_568_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX16 a_643_74_ a_363_74_ a_759_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX15 VDD GATE a_216_424_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX13 a_27_424_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX12 a_759_508_ a_817_48_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX9 a_363_74_ a_216_424_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 VDD a_817_48_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_817_48_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX0 a_568_392_ a_216_424_ a_643_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dllr_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dllr_1 D GATE_N Q Q_N RESET_B VDD VSS
*.PININFO D:B GATE_N:B Q:B Q_N:B RESET_B:B VDD:B VSS:B
MX19 VDD a_686_74_ a_889_92_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX17 a_802_508_ a_889_92_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX16 a_27_424_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX11 VDD a_27_424_ a_611_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX10 a_889_92_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 a_686_74_ a_231_74_ a_802_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX7 VDD GATE_N a_231_74_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX6 a_1437_112_ a_889_92_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 a_611_392_ a_373_74_ a_686_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX3 VDD a_889_92_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_373_74_ a_231_74_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 VDD a_1437_112_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX23 VSS a_1437_112_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 a_373_74_ a_231_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX21 a_889_92_ a_686_74_ a_1133_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
MX20 VSS GATE_N a_231_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 a_1437_112_ a_889_92_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX15 a_27_424_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX14 a_841_118_ a_889_92_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX13 VSS a_27_424_ a_608_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX12 a_686_74_ a_373_74_ a_841_118_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX8 VSS a_889_92_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_608_74_ a_231_74_ a_686_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX0 a_1133_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dllrq_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dllrq_1 D GATE_N Q RESET_B VDD VSS
*.PININFO D:B GATE_N:B Q:B RESET_B:B VDD:B VSS:B
MX18 a_357_392_ a_232_98_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 VSS a_897_406_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 a_654_392_ a_357_392_ a_854_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n 
+ ng=1
MX14 VSS a_27_136_ a_681_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX12 a_681_74_ a_232_98_ a_654_392_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n 
+ ng=1
MX9 a_27_136_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX6 a_1139_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_854_74_ a_897_406_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX3 a_897_406_ a_654_392_ a_1139_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n 
+ ng=1
MX1 VSS GATE_N a_232_98_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX19 VDD GATE_N a_232_98_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX15 a_897_406_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX13 a_654_392_ a_232_98_ a_793_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n 
+ ng=1
MX11 a_793_508_ a_897_406_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX10 VDD a_897_406_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX8 a_27_136_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 VDD a_27_136_ a_570_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 VDD a_654_392_ a_897_406_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX2 a_570_392_ a_357_392_ a_654_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n 
+ ng=1
MX0 a_357_392_ a_232_98_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_ebufn_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_ebufn_2 A TE_B VDD VSS Z
*.PININFO A:B TE_B:B VDD:B VSS:B Z:B
MX10 VSS A a_84_48_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 a_283_48_ TE_B VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX7 a_27_74_ a_84_48_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 a_27_74_ a_283_48_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 VSS a_283_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 Z a_84_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 VDD A a_84_48_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX9 VDD TE_B a_33_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX4 a_283_48_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX3 a_33_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Z a_84_48_ a_33_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX0 a_33_368_ a_84_48_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_ebufn_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_ebufn_4 A TE_B VDD VSS Z
*.PININFO A:B TE_B:B VDD:B VSS:B Z:B
MX19 a_378_74_ a_27_368_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 Z a_27_368_ a_378_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 a_378_74_ a_27_368_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX15 VSS a_208_74_ a_378_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX14 VSS TE_B a_208_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX13 a_378_74_ a_208_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 VSS a_208_74_ a_378_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 Z a_27_368_ a_378_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_27_368_ A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 a_378_74_ a_208_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 Z a_27_368_ a_348_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 a_348_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX10 Z a_27_368_ a_348_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 a_27_368_ A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX8 a_348_368_ a_27_368_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 a_348_368_ a_27_368_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 VDD TE_B a_208_74_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 a_348_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 VDD TE_B a_348_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX0 VDD TE_B a_348_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_ebufn_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_ebufn_8 A TE_B VDD VSS Z
*.PININFO A:B TE_B:B VDD:B VSS:B Z:B
MX0 a_28_368_ a_84_48_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 a_28_368_ a_84_48_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX13 Z a_84_48_ a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX18 a_28_368_ a_84_48_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX19 Z a_84_48_ a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX20 a_28_368_ a_84_48_ Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX27 Z a_84_48_ a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX33 Z a_84_48_ a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX37 a_833_48_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 a_84_48_ A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 VDD A a_84_48_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX8 a_28_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 VDD TE_B a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 a_28_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX16 a_28_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX17 VDD TE_B a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX23 VDD TE_B a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX35 a_28_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX36 VDD TE_B a_28_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Z a_84_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 Z a_84_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 Z a_84_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX24 a_27_74_ a_84_48_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX26 Z a_84_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX28 a_27_74_ a_84_48_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX32 a_27_74_ a_84_48_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX34 a_27_74_ a_84_48_ Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 VSS a_833_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 VSS a_833_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 a_27_74_ a_833_48_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX15 VSS a_833_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX21 a_27_74_ a_833_48_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX29 a_27_74_ a_833_48_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX30 a_27_74_ a_833_48_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX31 VSS a_833_48_ a_27_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX14 a_84_48_ A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX25 VSS A a_84_48_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 a_833_48_ TE_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_einvn_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_einvn_2 A TE_B VDD VSS Z
*.PININFO A:B TE_B:B VDD:B VSS:B Z:B
MX9 VSS TE_B a_115_464_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX6 Z A a_231_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_231_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS a_115_464_ a_231_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 a_231_74_ a_115_464_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 a_227_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 a_227_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX4 VDD TE_B a_115_464_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX1 VDD TE_B a_227_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX0 Z A a_227_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_einvn_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_einvn_4 A TE_B VDD VSS Z
*.PININFO A:B TE_B:B VDD:B VSS:B Z:B
MX17 VSS a_114_74_ a_281_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX15 a_281_74_ a_114_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX14 VSS TE_B a_114_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX13 a_281_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 VSS a_114_74_ a_281_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 Z A a_281_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 a_281_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 Z A a_281_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 a_281_74_ a_114_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 a_241_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 a_241_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX10 a_241_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 a_241_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 VDD TE_B a_241_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 VDD TE_B a_114_74_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX4 VDD TE_B a_241_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 Z A a_241_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX0 Z A a_241_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_einvn_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_einvn_8 A TE_B VDD VSS Z
*.PININFO A:B TE_B:B VDD:B VSS:B Z:B
MX0 Z A a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX14 Z A a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX16 a_239_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX18 a_239_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX26 a_239_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX27 Z A a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX29 a_239_368_ A Z VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX33 Z A a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX8 VDD TE_B a_126_74_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 a_239_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 VDD TE_B a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX13 a_239_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX20 VDD TE_B a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX23 a_239_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX24 a_239_368_ TE_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX25 VDD TE_B a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX30 VDD TE_B a_239_368_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_293_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 a_293_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 a_293_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 Z A a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 Z A a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX19 a_293_74_ A Z VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX21 Z A a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 Z A a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 VSS a_126_74_ a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_293_74_ a_126_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 a_293_74_ a_126_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX15 a_293_74_ a_126_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 VSS a_126_74_ a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX28 VSS a_126_74_ a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX31 a_293_74_ a_126_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX32 VSS a_126_74_ a_293_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS TE_B a_126_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_decap_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_decap_4 VDD VSS
*.PININFO VDD:B VSS:B
MX1 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
MX0 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_decap_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_decap_8 VDD VSS
*.PININFO VDD:B VSS:B
MX3 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
MX2 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
MX1 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
MX0 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_antennanp
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_antennanp A VDD VSS
*.PININFO A:I VDD:B VSS:B
Ddn_1 VSS A dantenna m=1 w=780n l=780n a=608.4f p=3.12u
DD0 A VDD dpantenna m=1 w=1.05u l=1.34u a=1.407p p=4.78u
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_tiehi
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_tiehi L_LO VDD VSS
*.PININFO L_LO:O VDD:B VSS:B
MMN2 net3 net2 VSS VSS sg13_lv_nmos m=1 w=795.00n l=130.00n ng=1
MMN1 net1 net1 VSS VSS sg13_lv_nmos m=1 w=300n l=130.00n ng=1
MMP2 L_LO net3 VDD VDD sg13_lv_pmos m=1 w=1.155u l=130.00n ng=1
MMP1 net2 net1 VDD VDD sg13_lv_pmos m=1 w=660.0n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_tielo
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_tielo L_LO VDD VSS
*.PININFO L_LO:O VDD:B VSS:B
MMN1 net3 net2 VSS VSS sg13_lv_nmos m=1 w=385.00n l=130.00n ng=1
MMN2 L_LO net1 VSS VSS sg13_lv_nmos m=1 w=880.0n l=130.00n ng=1
MMP1 net2 net2 VDD VDD sg13_lv_pmos m=1 w=300n l=130.00n ng=1
MMP2 net1 net3 VDD VDD sg13_lv_pmos m=1 w=1.045u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_sighold
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_sighold SIG VDD VSS
*.PININFO SIG:B VDD:B VSS:B
MN0 net1 SIG VSS VSS sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1
MN1 SIG net1 VSS VSS sg13_lv_nmos m=1 w=300.0n l=700.0n ng=1
MP0 net1 SIG VDD VDD sg13_lv_pmos m=1 w=450.00n l=130.00n ng=1
MP1 SIG net1 VDD VDD sg13_lv_pmos m=1 w=300.0n l=700.0n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_stdcell_allcells
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_stdcell_allcells
*.PININFO
XI1 net1 net2 VSS VDD net5 / sg13g2_and2_1
XI2 net6 net7 net8 VSS VDD net11 / sg13g2_and3_1
XI3 net12 net13 net14 net15 VSS VDD net18 / sg13g2_and4_1
XI4 net19 VDD VSS net20 / sg13g2_buf_1
XI5 net23 VDD VSS net24 / sg13g2_buf_16
XI6 net27 VDD VSS net28 / sg13g2_buf_2
XI7 net31 VDD VSS net32 / sg13g2_buf_4
XI8 net35 VDD VSS net36 / sg13g2_buf_8
XI9 net39 net40 net41 VSS VDD net44 net45 / sg13g2_dfrbp_2
XI10 net46 VSS VDD net49 / sg13g2_dlygate4sd1_1
XI11 net50 VSS VDD net53 / sg13g2_dlygate4sd2_1
XI12 net54 VSS VDD net57 / sg13g2_dlygate4sd3_1
XI13 net61 VDD VSS net58 / sg13g2_inv_1
XI14 net62 VSS VDD net65 / sg13g2_inv_16
XI15 net66 VDD VSS net69 / sg13g2_inv_2
XI16 net70 VSS VDD net73 / sg13g2_inv_4
XI17 net74 VSS VDD net77 / sg13g2_inv_8
XI18 net78 net79 net80 VSS VDD net83 / sg13g2_mux2_1
XI19 net84 net85 net86 VSS VDD net89 / sg13g2_a21o_1
XI20 net90 net91 net92 net93 net94 net95 VSS VDD net98 / sg13g2_mux4_1
XI21 net99 net100 VSS VDD net103 / sg13g2_nand2_1
XI22 net104 net105 VSS VDD net108 / sg13g2_nand2b_1
XI23 net109 net110 net111 VSS VDD net114 / sg13g2_nand3b_1
XI24 net115 net116 VSS VDD net119 / sg13g2_nor2_1
XI25 net120 net121 net122 VSS VDD net125 / sg13g2_nor3_1
XI26 net126 net127 net128 net129 VSS VDD net132 / sg13g2_nor4_1
XI27 net133 net134 VDD VSS net137 / sg13g2_or2_1
XI28 net138 net139 net140 VSS VDD net143 / sg13g2_or3_1
XI29 net147 net146 net145 net144 VDD VSS net148 / sg13g2_or4_1
XI30 net151 net152 VSS VDD net155 / sg13g2_xnor2_1
XI31 net156 net157 VSS VDD net160 / sg13g2_xor2_1
XI32 net161 net162 net166 net167 net163 VDD VSS / sg13g2_dfrbp_1
XI33 net168 net169 net176 net177 net170 net171 net172 net173 VDD VSS / 
+ sg13g2_sdfbbp_1
XI34 net178 net179 net182 VDD VSS / sg13g2_lgcp_1
XI35 net183 net184 net186 net185 VDD VSS / sg13g2_slgcp_1
XI36 net189 net190 net193 VDD VSS / sg13g2_dlhq_1
XI37 net194 net195 net199 net200 net196 VDD VSS / sg13g2_dlhr_1
XI38 net201 net202 net206 net203 VDD VSS / sg13g2_dlhrq_1
XI39 net207 net208 net212 net213 net209 VDD VSS / sg13g2_dllr_1
XI40 net214 net215 net219 net216 VDD VSS / sg13g2_dllrq_1
XI41 net220 net221 VDD VSS net224 / sg13g2_ebufn_2
XI42 net225 net226 VDD VSS net229 / sg13g2_ebufn_4
XI43 net230 net231 VDD VSS net234 / sg13g2_ebufn_8
XI44 net235 net236 VDD VSS net239 / sg13g2_einvn_2
XI45 net240 net241 VDD VSS net244 / sg13g2_einvn_4
XI46 net245 net246 VDD VSS net249 / sg13g2_einvn_8
XI0 VDD VSS / sg13g2_decap_4
XI47 VDD VSS / sg13g2_decap_8
XI48 net3 VDD VSS / sg13g2_antennanp
XI49 net4 VDD VSS / sg13g2_tiehi
XI50 net9 VDD VSS / sg13g2_tielo
XI51 net10 VDD VSS / sg13g2_sighold
.ENDS

