########################################################################
#
# Copyright 2023 IHP PDK Authors
# 
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
# 
#    https://www.apache.org/licenses/LICENSE-2.0
# 
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
########################################################################

VERSION 5.7 ;
BUSBITCHARS "<>" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SIZE        0.48 BY 3.78 ;
END  CoreSite

MACRO sg13g2_a21o_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21o_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.81 0.405 3.215 0.965 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.215 1.565 2.545 2 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.57 2.005 2 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6159 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.885 1.225 1.145 ;
        RECT 0.205 2.095 0.56 3.105 ;
        RECT 0.205 0.885 0.445 3.105 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.405 2.585 2.665 4 ;
        RECT 0.81 2.14 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.92 1.145 3.165 1.41 ;
        RECT 2.455 1.145 3.165 1.31 ;
        RECT 2.455 -0.22 2.615 1.31 ;
        RECT 1.455 -0.22 1.715 0.965 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.915 2.21 3.175 3.125 ;
      RECT 1.855 2.21 2.115 3.125 ;
      RECT 1.855 2.21 3.175 2.405 ;
      RECT 1.335 2.17 1.595 3.125 ;
      RECT 1.335 1.54 1.575 3.125 ;
      RECT 1.415 1.22 1.575 3.125 ;
      RECT 0.625 1.54 1.575 1.87 ;
      RECT 1.415 1.22 2.27 1.385 ;
      RECT 2.02 0.825 2.27 1.385 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21o_1

MACRO sg13g2_a21o_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21o_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.2 1.565 3.69 2 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.69 1.565 3.02 2 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.23 1.57 2.48 2 ;
    END
  END B1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 0.74 1.045 3.16 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.88 2.585 3.14 4 ;
        RECT 1.295 2.18 1.555 4 ;
        RECT 0.275 2.18 0.535 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.4 -0.22 3.645 1.385 ;
        RECT 1.935 -0.22 2.195 0.99 ;
        RECT 1.295 -0.22 1.555 1.37 ;
        RECT 0.275 -0.22 0.535 1.37 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 3.39 2.21 3.65 3.125 ;
      RECT 2.33 2.21 2.59 3.125 ;
      RECT 2.33 2.21 3.65 2.405 ;
      RECT 1.81 2.17 2.07 3.125 ;
      RECT 1.81 1.22 2.05 3.125 ;
      RECT 1.235 1.67 2.05 1.93 ;
      RECT 1.81 1.22 2.745 1.385 ;
      RECT 2.495 0.725 2.745 1.385 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21o_2

MACRO sg13g2_a21oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21oi_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.835 -0.22 2.095 1.37 ;
        RECT 0.305 -0.22 0.565 0.93 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.325 2.9 1.585 4 ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.07 1.62 1.585 1.83 ;
        RECT 1.325 0.77 1.585 1.83 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.55 2.095 1.95 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 0.77 1.075 1.37 ;
        RECT 0.305 2.13 0.89 2.29 ;
        RECT 0.715 1.21 0.89 2.29 ;
        RECT 0.305 2.13 0.565 3.11 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.155 0.53 1.9 ;
    END
  END B1
  OBS
    LAYER Metal1 ;
      RECT 1.835 2.13 2.095 3.11 ;
      RECT 0.815 2.555 1.075 3.11 ;
      RECT 1.075 2.13 2.095 2.715 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21oi_1

MACRO sg13g2_a21oi_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a21oi_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.315 -0.22 3.575 1.42 ;
        RECT 2.295 -0.22 2.555 0.98 ;
        RECT 0.255 -0.22 0.515 1.42 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 1.785 2.95 2.045 4 ;
        RECT 0.765 2.95 1.025 4 ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.28 1.625 3.575 2.28 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.988 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.805 0.72 3.065 2.715 ;
        RECT 1.275 1.16 3.065 1.39 ;
        RECT 1.275 0.85 1.535 1.39 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 2.09 2.3 2.315 ;
        RECT 2.04 1.6 2.3 2.315 ;
        RECT 0.39 1.6 0.77 2.315 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 1.57 1.725 1.9 ;
    END
  END A1
  OBS
    LAYER Metal1 ;
      RECT 2.295 2.9 3.575 3.16 ;
      RECT 3.315 2.505 3.575 3.16 ;
      RECT 1.275 2.505 1.535 3.16 ;
      RECT 0.255 2.505 0.515 3.16 ;
      RECT 2.295 2.505 2.555 3.16 ;
      RECT 0.255 2.505 2.555 2.765 ;
      RECT 1.785 0.445 2.045 0.98 ;
      RECT 0.765 0.445 1.025 0.98 ;
      RECT 0.765 0.445 2.045 0.67 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a21oi_2

MACRO sg13g2_a221oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a221oi_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.32 -0.22 3.58 0.98 ;
        RECT 0.77 -0.22 1.03 0.98 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.32 2.505 3.58 4 ;
        RECT 2.3 2.9 2.56 4 ;
    END
  END VDD
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.88 1.57 1.36 1.9 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 1.57 0.64 1.9 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.54 1.57 2 1.9 ;
        RECT 1.72 1.16 2 1.9 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.18 1.57 2.7 1.9 ;
        RECT 2.18 1.16 2.48 1.9 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1356 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 2.08 3.745 2.29 ;
        RECT 3.565 1.16 3.745 2.29 ;
        RECT 2.81 1.16 3.745 1.37 ;
        RECT 2.81 0.72 3.07 1.37 ;
        RECT 1.28 0.72 3.07 0.98 ;
        RECT 0.26 1.16 1.54 1.37 ;
        RECT 1.28 0.72 1.54 1.37 ;
        RECT 0.26 2.08 0.52 3.16 ;
        RECT 0.26 0.72 0.52 1.37 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.88 1.57 3.385 1.9 ;
    END
  END A2
  OBS
    LAYER Metal1 ;
      RECT 2.81 2.505 3.07 3.16 ;
      RECT 1.28 2.505 1.54 2.765 ;
      RECT 1.28 2.505 3.07 2.715 ;
      RECT 0.77 2.95 2.05 3.16 ;
      RECT 1.79 2.9 2.05 3.16 ;
      RECT 0.77 2.505 1.03 3.16 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a221oi_1

MACRO sg13g2_a22oi_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_a22oi_1 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9584 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 0.89 1.75 1.15 ;
        RECT 1.31 2.25 1.6 2.9 ;
        RECT 1.42 0.89 1.6 2.9 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 1.33 1.24 2.07 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 1.7 2.08 2.44 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.42 1.33 2.72 2.07 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 1.36 2.09 1.52 ;
        RECT 1.93 0.55 2.09 1.52 ;
        RECT 0.62 0.55 2.09 0.71 ;
        RECT 0.17 1.33 0.78 1.49 ;
        RECT 0.62 0.55 0.78 1.49 ;
        RECT 0.17 1.33 0.47 2.07 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.44 2.25 2.7 4 ;
        RECT 0.18 2.25 0.45 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.44 -0.22 2.7 1.15 ;
        RECT 0.18 -0.22 0.44 1.15 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.8 3.085 2.08 3.33 ;
      RECT 1.82 2.62 2.08 3.33 ;
      RECT 0.8 2.25 1.06 3.33 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_a22oi_1

MACRO sg13g2_and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and2_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.105 0.405 0.78 0.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 1.435 1.17 1.87 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.775 2.14 2.275 3.11 ;
        RECT 2.04 0.78 2.275 3.11 ;
        RECT 1.775 0.78 2.275 1.36 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.265 2.485 1.525 4 ;
        RECT 0.245 2.425 0.505 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.265 -0.22 1.525 1.155 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.755 2.05 1.015 3.11 ;
      RECT 0.245 2.05 1.56 2.24 ;
      RECT 1.4 1.57 1.56 2.24 ;
      RECT 0.245 1.14 0.505 2.24 ;
      RECT 1.4 1.57 1.74 1.9 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and2_1

MACRO sg13g2_and2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.105 0.405 0.78 0.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 1.435 1.17 1.87 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.775 2.14 2.105 3.11 ;
        RECT 1.92 0.78 2.105 3.11 ;
        RECT 1.775 0.78 2.105 1.36 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.285 2.485 2.545 4 ;
        RECT 1.265 2.485 1.525 4 ;
        RECT 0.245 2.425 0.505 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.285 -0.22 2.545 1.155 ;
        RECT 1.265 -0.22 1.525 1.155 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.755 2.05 1.015 3.11 ;
      RECT 0.245 2.05 1.56 2.24 ;
      RECT 1.4 1.57 1.56 2.24 ;
      RECT 0.245 1.14 0.505 2.24 ;
      RECT 1.4 1.57 1.74 1.9 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and2_2

MACRO sg13g2_and3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and3_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.78 2.17 3.065 3.27 ;
        RECT 2.895 1.125 3.065 3.27 ;
        RECT 2.44 1.125 3.065 1.385 ;
        RECT 2.44 0.77 2.7 1.385 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 0.475 1.59 1.09 ;
        RECT 0.35 0.475 1.59 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.4 1.54 1.98 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 1.4 2.06 1.95 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 1.93 2.615 2.53 4 ;
        RECT 0.91 2.73 1.17 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 1.93 -0.22 2.19 1.14 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.4 1.09 0.66 3.115 ;
      RECT 1.42 2.16 1.68 3.085 ;
      RECT 0.4 2.16 2.405 2.32 ;
      RECT 2.245 1.57 2.405 2.32 ;
      RECT 2.245 1.57 2.645 1.9 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and3_1

MACRO sg13g2_and3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and3_2 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 2.51 3.065 2.69 ;
        RECT 2.835 1.29 3.065 2.69 ;
        RECT 2.44 1.29 3.065 1.55 ;
        RECT 2.435 2.51 2.705 3.36 ;
        RECT 2.44 0.77 2.7 1.55 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 0.475 1.59 1.09 ;
        RECT 0.35 0.475 1.59 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.4 1.54 1.98 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 1.4 2.06 1.95 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.955 2.875 3.225 4 ;
        RECT 1.93 2.615 2.19 4 ;
        RECT 0.91 2.73 1.17 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.95 -0.22 3.21 1.09 ;
        RECT 1.93 -0.22 2.19 1.14 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.4 1.09 0.66 3.115 ;
      RECT 1.42 2.16 1.68 3.085 ;
      RECT 0.4 2.16 2.405 2.32 ;
      RECT 2.245 1.735 2.405 2.32 ;
      RECT 2.245 1.735 2.645 2.065 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and3_2

MACRO sg13g2_and4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and4_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.35 1.07 2.01 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 0.66 1.565 2.025 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.66 2.125 2.01 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 1.57 2.665 2 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8928 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 2.07 3.685 3.12 ;
        RECT 3.525 0.64 3.685 3.12 ;
        RECT 3.205 0.64 3.685 1.26 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.54 2.585 2.8 4 ;
        RECT 1.445 2.56 1.705 4 ;
        RECT 0.425 2.56 0.685 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.55 -0.22 2.815 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.935 2.22 1.195 3.125 ;
      RECT 1.985 2.22 2.245 3.12 ;
      RECT 0.355 2.22 3.01 2.38 ;
      RECT 2.85 1.54 3.01 2.38 ;
      RECT 0.355 0.645 0.525 2.38 ;
      RECT 2.85 1.54 3.205 1.87 ;
      RECT 0.355 0.645 0.995 1.17 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and4_1

MACRO sg13g2_and4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_and4_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.35 1.07 2.01 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 0.66 1.565 2.025 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.66 2.125 2.01 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 1.57 2.665 2 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9672 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 2.07 3.685 3.12 ;
        RECT 3.525 0.64 3.685 3.12 ;
        RECT 3.205 0.64 3.685 1.26 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 3.865 2.13 4.125 4 ;
        RECT 2.54 2.585 2.8 4 ;
        RECT 1.445 2.56 1.705 4 ;
        RECT 0.425 2.56 0.685 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 3.865 -0.22 4.125 1.26 ;
        RECT 2.55 -0.22 2.815 1.21 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.935 2.22 1.195 3.125 ;
      RECT 1.985 2.22 2.245 3.12 ;
      RECT 0.355 2.22 3.01 2.38 ;
      RECT 2.85 1.54 3.01 2.38 ;
      RECT 0.355 0.645 0.525 2.38 ;
      RECT 2.85 1.54 3.205 1.87 ;
      RECT 0.355 0.645 0.995 1.17 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_and4_2

MACRO sg13g2_antennanp
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_antennanp 0 0 ;
  SIZE 1.44 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.44 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.44 0.22 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0154 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.57 1.05 1.16 ;
        RECT 0.38 1.13 0.63 2.41 ;
    END
  END A
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_antennanp

MACRO sg13g2_buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_1 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.1 1.65 0.87 2.115 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6548 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.49 2.02 1.79 3.18 ;
        RECT 1.6 0.55 1.79 3.18 ;
        RECT 1.5 0.55 1.79 1.29 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.945 2.84 1.245 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.935 -0.22 1.265 1.025 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.43 2.44 0.7 3.18 ;
      RECT 0.43 2.44 1.26 2.62 ;
      RECT 1.09 1.29 1.26 2.62 ;
      RECT 1.09 1.5 1.415 1.83 ;
      RECT 0.315 1.29 1.26 1.465 ;
      RECT 0.315 1 0.705 1.465 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_1

MACRO sg13g2_buf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_16 0 0 ;
  SIZE 12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    ANTENNADIFFAREA 5.6544 LAYER Metal2 ;
    PORT
      LAYER Metal1 ;
        RECT 7.91 0.64 8.17 3.105 ;
        RECT 6.89 0.645 7.15 3.105 ;
        RECT 5.87 0.65 6.13 3.105 ;
        RECT 4.85 0.635 5.11 3.11 ;
        RECT 3.83 0.65 4.09 3.11 ;
        RECT 2.81 0.645 3.07 3.11 ;
        RECT 1.79 0.645 2.05 3.11 ;
        RECT 0.77 0.64 1.03 3.105 ;
      LAYER Metal2 ;
        RECT 0.745 2.405 8.195 2.635 ;
      LAYER Via1 ;
        RECT 0.805 2.425 0.995 2.615 ;
        RECT 1.825 2.425 2.015 2.615 ;
        RECT 2.845 2.425 3.035 2.615 ;
        RECT 3.865 2.425 4.055 2.615 ;
        RECT 4.885 2.425 5.075 2.615 ;
        RECT 5.91 2.425 6.1 2.615 ;
        RECT 6.925 2.425 7.115 2.615 ;
        RECT 7.95 2.425 8.14 2.615 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.4508 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.78 1.57 11.44 1.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 12 4 ;
        RECT 11.48 2.205 11.74 4 ;
        RECT 10.46 2.545 10.72 4 ;
        RECT 9.44 2.54 9.7 4 ;
        RECT 8.42 2.54 8.68 4 ;
        RECT 7.4 2.145 7.66 4 ;
        RECT 6.38 2.145 6.64 4 ;
        RECT 5.36 2.145 5.62 4 ;
        RECT 4.34 2.145 4.6 4 ;
        RECT 3.32 2.14 3.58 4 ;
        RECT 2.3 2.14 2.56 4 ;
        RECT 1.28 2.14 1.54 4 ;
        RECT 0.26 2.14 0.52 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 12 0.22 ;
        RECT 11.48 -0.22 11.74 1.235 ;
        RECT 10.46 -0.22 10.72 0.995 ;
        RECT 9.44 -0.22 9.7 1 ;
        RECT 8.42 -0.22 8.685 0.99 ;
        RECT 7.4 -0.22 7.66 1.28 ;
        RECT 6.38 -0.22 6.64 1.18 ;
        RECT 5.36 -0.22 5.62 1.275 ;
        RECT 4.34 -0.22 4.6 1.27 ;
        RECT 3.32 -0.22 3.58 1.195 ;
        RECT 2.3 -0.22 2.56 1.275 ;
        RECT 1.28 -0.22 1.54 1.28 ;
        RECT 0.26 -0.22 0.52 1.27 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 10.97 2.17 11.23 3.105 ;
      RECT 9.95 2.17 10.21 3.105 ;
      RECT 8.93 2.17 9.19 3.105 ;
      RECT 8.385 2.17 11.23 2.34 ;
      RECT 8.385 1.18 8.595 2.34 ;
      RECT 8.385 1.18 11.23 1.35 ;
      RECT 10.97 0.645 11.23 1.35 ;
      RECT 9.95 0.64 10.21 1.35 ;
      RECT 8.93 0.645 9.19 1.35 ;
      RECT 7.38 1.52 7.665 1.95 ;
      RECT 6.37 1.52 6.655 1.95 ;
      RECT 5.335 1.52 5.62 1.95 ;
      RECT 4.33 1.52 4.615 1.95 ;
      RECT 3.3 1.52 3.595 1.95 ;
      RECT 2.28 1.52 2.565 1.95 ;
      RECT 1.24 1.52 1.55 1.955 ;
    LAYER Via1 ;
      RECT 8.395 1.59 8.585 1.78 ;
      RECT 7.435 1.59 7.625 1.78 ;
      RECT 6.415 1.59 6.605 1.78 ;
      RECT 5.395 1.59 5.585 1.78 ;
      RECT 4.375 1.59 4.565 1.78 ;
      RECT 3.355 1.59 3.545 1.78 ;
      RECT 2.335 1.59 2.525 1.78 ;
      RECT 1.315 1.59 1.505 1.78 ;
    LAYER Metal2 ;
      RECT 1.24 1.57 8.645 1.8 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_16

MACRO sg13g2_buf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_2 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 1.57 2.275 2 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.945 0.635 1.275 2.37 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.485 2.895 1.745 4 ;
        RECT 0.15 2.12 0.41 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.485 -0.22 1.745 0.995 ;
        RECT 0.465 -0.22 0.725 1.275 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.97 2.18 2.26 3.1 ;
      RECT 0.605 2.55 2.26 2.71 ;
      RECT 1.495 1.23 1.655 2.71 ;
      RECT 0.605 1.52 0.765 2.71 ;
      RECT 0.105 1.52 0.765 1.85 ;
      RECT 1.495 1.23 2.255 1.39 ;
      RECT 1.995 0.72 2.255 1.39 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_2

MACRO sg13g2_buf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_4 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.995 2.025 3.13 ;
        RECT 0.745 1.065 2.025 1.285 ;
        RECT 1.765 0.645 2.025 1.285 ;
        RECT 0.745 1.995 2.025 2.165 ;
        RECT 0.745 0.63 1.005 3.13 ;
    END
  END X
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.77 1.57 3.15 2 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.295 2.64 3.555 4 ;
        RECT 2.275 2.285 2.535 4 ;
        RECT 1.255 2.345 1.515 4 ;
        RECT 0.235 2.115 0.495 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.41 0.595 2.94 0.87 ;
        RECT 2.545 -0.22 2.805 0.87 ;
        RECT 1.255 -0.22 1.515 0.88 ;
        RECT 0.235 -0.22 0.495 1 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.785 2.205 3.045 2.77 ;
      RECT 2.785 2.205 3.59 2.42 ;
      RECT 3.4 0.64 3.59 2.42 ;
      RECT 1.305 1.555 2.53 1.815 ;
      RECT 2.36 1.18 2.53 1.815 ;
      RECT 2.36 1.18 3.59 1.35 ;
      RECT 3.245 0.64 3.59 1.35 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_4

MACRO sg13g2_buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_buf_8 0 0 ;
  SIZE 6.24 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.7254 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 1.57 1.55 1.95 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8272 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.65 5.52 3.12 ;
        RECT 2.2 2.07 5.52 2.23 ;
        RECT 2.2 1.13 5.52 1.3 ;
        RECT 4.24 2.07 4.5 3.13 ;
        RECT 4.24 0.645 4.5 1.3 ;
        RECT 3.22 2.07 3.48 3.125 ;
        RECT 3.22 0.64 3.48 1.3 ;
        RECT 2.2 2.07 2.46 3.12 ;
        RECT 2.2 0.645 2.46 1.3 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 6.24 4 ;
        RECT 5.77 2.12 6.03 4 ;
        RECT 4.75 2.42 5.01 4 ;
        RECT 3.73 2.43 3.99 4 ;
        RECT 2.71 2.43 2.97 4 ;
        RECT 1.69 2.575 1.95 4 ;
        RECT 0.67 2.575 0.93 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 6.24 0.22 ;
        RECT 5.77 -0.22 6.03 1.275 ;
        RECT 4.75 -0.22 5.01 0.945 ;
        RECT 3.73 -0.22 3.99 0.95 ;
        RECT 2.71 -0.22 2.97 0.95 ;
        RECT 1.69 -0.22 1.95 0.99 ;
        RECT 0.67 -0.22 0.93 0.995 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.18 2.17 1.44 3.125 ;
      RECT 0.16 2.17 0.42 3.125 ;
      RECT 0.16 2.17 1.94 2.34 ;
      RECT 1.77 1.18 1.94 2.34 ;
      RECT 1.77 1.555 4.975 1.815 ;
      RECT 0.16 1.18 1.94 1.35 ;
      RECT 1.18 0.645 1.44 1.35 ;
      RECT 0.16 0.64 0.42 1.35 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_buf_8

MACRO sg13g2_decap_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_decap_4 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 1.065 2.54 1.79 4 ;
        RECT 1.065 1.47 1.405 4 ;
        RECT 0.13 2.535 0.4 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 1.51 -0.22 1.79 0.935 ;
        RECT 0.53 -0.22 0.855 1.805 ;
        RECT 0.13 -0.22 0.855 0.935 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_decap_4

MACRO sg13g2_decap_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_decap_8 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.945 2.21 3.205 4 ;
        RECT 1.22 1.475 2.155 4 ;
        RECT 0.185 2.205 0.445 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.585 -0.22 3.195 0.99 ;
        RECT 2.585 -0.22 2.835 1.81 ;
        RECT 1.53 -0.22 1.835 1.03 ;
        RECT 0.52 -0.22 0.81 1.81 ;
        RECT 0.175 -0.22 0.81 0.99 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_decap_8

MACRO sg13g2_dfrbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dfrbp_1 0 0 ;
  SIZE 12.48 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 1.575 2.49 1.985 ;
        RECT 2.045 1.575 2.49 1.915 ;
    END
  END CLK
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal2 ;
      ANTENNAMAXAREACAR 1.208791 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.330586 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.325 2.055 8.725 2.385 ;
        RECT 5.615 2.045 6.015 2.355 ;
        RECT 1.255 1.35 1.525 2.36 ;
      LAYER Metal2 ;
        RECT 8.275 2 8.725 2.37 ;
        RECT 1.28 2 8.725 2.2 ;
        RECT 5.6 2 5.89 2.37 ;
        RECT 1.28 1.965 1.57 2.37 ;
      LAYER Via1 ;
        RECT 1.305 2.015 1.495 2.205 ;
        RECT 5.665 2.13 5.855 2.32 ;
        RECT 8.44 2.145 8.63 2.335 ;
    END
  END RESET_B
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 1.22 0.735 2.415 ;
    END
  END D
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0391 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.79 2.08 10.38 3.165 ;
        RECT 10.09 0.605 10.35 3.165 ;
    END
  END Q_N
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.785 2.08 12.145 3.16 ;
        RECT 11.975 0.645 12.145 3.16 ;
        RECT 11.775 0.645 12.145 1.28 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 12.48 4 ;
        RECT 11.255 2.52 11.515 4 ;
        RECT 9.25 2.395 9.51 4 ;
        RECT 8.245 2.65 8.415 4 ;
        RECT 6.235 1.99 6.415 4 ;
        RECT 4.98 2.875 5.24 4 ;
        RECT 2.395 2.94 2.655 4 ;
        RECT 1.375 2.935 1.635 4 ;
        RECT 0.355 2.86 0.615 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 12.48 0.22 ;
        RECT 11.285 -0.22 11.545 1.27 ;
        RECT 9.545 -0.22 9.805 0.86 ;
        RECT 8.13 -0.22 8.39 0.875 ;
        RECT 5.48 -0.22 5.74 0.63 ;
        RECT 2.425 -0.22 2.685 1.02 ;
        RECT 1.28 -0.22 1.54 0.91 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 10.745 0.705 11.005 3.135 ;
      RECT 10.745 1.52 11.77 1.85 ;
      RECT 10.745 0.705 11.01 1.85 ;
      RECT 8.71 2.645 9.065 2.91 ;
      RECT 8.905 1.995 9.065 2.91 ;
      RECT 8.905 1.995 9.6 2.155 ;
      RECT 9.435 1.12 9.6 2.155 ;
      RECT 7.96 1.12 8.22 1.375 ;
      RECT 7.96 1.12 9.6 1.29 ;
      RECT 9.015 0.665 9.275 1.29 ;
      RECT 7.255 2.615 8.065 2.875 ;
      RECT 7.905 1.645 8.065 2.875 ;
      RECT 7.6 1.645 9.12 1.815 ;
      RECT 8.85 1.5 9.12 1.815 ;
      RECT 7.6 0.67 7.77 1.815 ;
      RECT 7.16 0.67 7.77 0.885 ;
      RECT 7.14 2.085 7.725 2.415 ;
      RECT 2.905 2.085 3.165 2.415 ;
      RECT 2.905 2.085 3.225 2.3 ;
      RECT 2.905 2.085 3.245 2.285 ;
      RECT 2.905 2.085 3.25 2.28 ;
      RECT 2.905 2.085 3.275 2.26 ;
      RECT 2.905 2.085 3.515 2.215 ;
      RECT 3.37 1.875 4 2.17 ;
      RECT 7.14 1.12 7.3 2.415 ;
      RECT 3.14 2.045 4 2.17 ;
      RECT 3.37 1.31 3.53 2.17 ;
      RECT 3.25 0.475 3.415 1.47 ;
      RECT 6.795 1.12 7.3 1.45 ;
      RECT 6.795 0.53 6.965 1.45 ;
      RECT 2.92 0.765 3.415 1.055 ;
      RECT 5.005 0.81 6.08 0.97 ;
      RECT 5.92 0.53 6.08 0.97 ;
      RECT 5.005 0.475 5.19 0.97 ;
      RECT 5.92 0.53 6.965 0.695 ;
      RECT 3.25 0.475 5.19 0.635 ;
      RECT 6.745 1.63 6.925 2.935 ;
      RECT 4.86 1.15 5.095 2.345 ;
      RECT 6.215 1.63 6.925 1.79 ;
      RECT 6.215 1.15 6.48 1.79 ;
      RECT 6.265 0.88 6.48 1.79 ;
      RECT 4.86 1.15 6.48 1.31 ;
      RECT 4.045 2.7 4.68 2.915 ;
      RECT 4.52 0.89 4.68 2.915 ;
      RECT 5.525 2.535 5.785 2.86 ;
      RECT 4.52 2.535 5.785 2.695 ;
      RECT 5.275 1.665 5.435 2.695 ;
      RECT 5.275 1.665 6.03 1.835 ;
      RECT 5.74 1.505 6.03 1.835 ;
      RECT 4.195 0.89 4.68 1.175 ;
      RECT 0.865 2.625 1.125 3.095 ;
      RECT 3.555 2.595 3.82 2.91 ;
      RECT 3.63 2.36 3.82 2.91 ;
      RECT 0.915 2.595 3.82 2.755 ;
      RECT 0.915 0.76 1.075 3.095 ;
      RECT 3.63 2.36 4.34 2.52 ;
      RECT 4.18 1.355 4.34 2.52 ;
      RECT 3.765 1.355 4.34 1.515 ;
      RECT 3.765 0.895 3.96 1.515 ;
      RECT 3.68 0.895 3.96 1.155 ;
      RECT 0.4 0.76 1.075 0.95 ;
      RECT 0.4 0.685 0.66 0.95 ;
      RECT 1.885 2.12 2.145 2.41 ;
      RECT 1.705 2.12 2.145 2.315 ;
      RECT 1.705 1.02 1.865 2.315 ;
      RECT 2.835 1.645 3.19 1.865 ;
      RECT 2.835 1.235 3.01 1.865 ;
      RECT 1.705 1.235 3.01 1.395 ;
      RECT 1.775 0.815 2.145 1.395 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dfrbp_1

MACRO sg13g2_dfrbp_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dfrbp_2 0 0 ;
  SIZE 14.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
      ANTENNAGATEAREA 0.3276 LAYER Metal2 ;
      ANTENNAMAXAREACAR 1.142857 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.330586 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.595 1.65 9.985 1.97 ;
        RECT 2.385 1.61 2.755 1.955 ;
        RECT 1.025 1.45 1.315 1.98 ;
      LAYER Metal2 ;
        RECT 1.075 2 9.93 2.2 ;
        RECT 9.64 1.735 9.93 2.2 ;
        RECT 2.43 1.705 2.72 2.2 ;
        RECT 1.075 1.58 1.275 2.2 ;
      LAYER Via1 ;
        RECT 1.08 1.66 1.27 1.85 ;
        RECT 2.48 1.755 2.67 1.945 ;
        RECT 9.69 1.77 9.88 1.96 ;
    END
  END RESET_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 14.4 0.22 ;
        RECT 13.935 -0.22 14.21 1.295 ;
        RECT 12.93 -0.22 13.19 1.29 ;
        RECT 11.91 -0.22 12.17 0.81 ;
        RECT 10.91 -0.22 11.155 1.27 ;
        RECT 9.51 -0.22 9.77 0.885 ;
        RECT 5.635 -0.22 5.91 0.66 ;
        RECT 2.345 -0.22 2.515 0.97 ;
        RECT 1.14 -0.22 1.41 0.975 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 14.4 4 ;
        RECT 13.59 2.06 13.84 4 ;
        RECT 12.56 2.07 12.815 4 ;
        RECT 11.465 1.975 11.725 4 ;
        RECT 10.45 2.495 10.725 4 ;
        RECT 9.33 2.505 9.595 4 ;
        RECT 6.16 2.955 6.445 4 ;
        RECT 2.945 2.86 3.115 4 ;
        RECT 0.15 2.215 0.46 4 ;
    END
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 1.07 0.5 1.77 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7124 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.19 1.515 13.72 1.775 ;
        RECT 13.42 0.545 13.72 1.775 ;
        RECT 13.07 2.04 13.36 3.175 ;
        RECT 13.19 1.515 13.36 3.175 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.395 0.99 11.93 1.61 ;
        RECT 11 1.52 11.78 1.74 ;
        RECT 11.395 0.55 11.66 1.74 ;
        RECT 11 1.52 11.19 3.1 ;
    END
  END Q_N
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal2 ;
      ANTENNAMAXAREACAR 0.508892 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.149297 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.76 1.335 6.99 1.87 ;
      LAYER Metal2 ;
        RECT 6.65 1.24 7.12 1.745 ;
      LAYER Via1 ;
        RECT 6.78 1.515 6.97 1.705 ;
    END
  END CLK
  OBS
    LAYER Metal1 ;
      RECT 11.95 1.94 12.36 2.98 ;
      RECT 12.19 1.355 12.36 2.98 ;
      RECT 12.19 1.515 13 1.83 ;
      RECT 12.19 1.355 12.685 1.83 ;
      RECT 12.4 0.55 12.685 1.83 ;
      RECT 9.935 2.15 10.14 2.555 ;
      RECT 9.13 2.15 10.14 2.32 ;
      RECT 9.13 2.15 10.73 2.31 ;
      RECT 10.57 0.55 10.73 2.31 ;
      RECT 9.13 1.655 9.385 2.32 ;
      RECT 10.26 0.55 10.73 0.945 ;
      RECT 8.455 2.125 8.66 2.5 ;
      RECT 8.455 2.125 8.95 2.295 ;
      RECT 8.79 1.145 8.95 2.295 ;
      RECT 10.165 1.275 10.39 1.625 ;
      RECT 8.79 1.275 10.39 1.465 ;
      RECT 7.96 1.145 8.97 1.315 ;
      RECT 7.51 0.805 7.68 1.31 ;
      RECT 7.51 0.805 9.29 0.965 ;
      RECT 9.04 0.55 9.29 0.965 ;
      RECT 7.745 1.555 7.935 2.925 ;
      RECT 1.495 2.485 1.97 2.655 ;
      RECT 1.495 1.215 1.655 2.655 ;
      RECT 2.935 1.755 3.23 1.965 ;
      RECT 2.935 1.215 3.095 1.965 ;
      RECT 7.17 1.555 7.935 1.725 ;
      RECT 7.17 0.465 7.33 1.725 ;
      RECT 1.495 1.215 3.095 1.385 ;
      RECT 2.705 0.485 2.875 1.385 ;
      RECT 1.655 0.815 1.975 1.385 ;
      RECT 5.295 0.84 6.255 1 ;
      RECT 6.09 0.465 6.255 1 ;
      RECT 5.295 0.485 5.455 1 ;
      RECT 2.705 0.485 5.455 0.645 ;
      RECT 6.09 0.465 8.82 0.625 ;
      RECT 7.315 3.105 8.275 3.265 ;
      RECT 8.115 1.5 8.275 3.265 ;
      RECT 5.425 2.06 5.785 3.18 ;
      RECT 7.315 2.59 7.505 3.265 ;
      RECT 5.425 2.59 7.505 2.77 ;
      RECT 4.72 2.11 5.785 2.44 ;
      RECT 5.145 2.06 5.785 2.44 ;
      RECT 5.145 1.18 5.42 2.44 ;
      RECT 8.115 1.5 8.605 1.805 ;
      RECT 6.15 2.055 7.56 2.37 ;
      RECT 6.15 1.54 6.32 2.37 ;
      RECT 5.65 1.54 6.32 1.87 ;
      RECT 5.65 1.54 6.58 1.845 ;
      RECT 6.42 1.075 6.58 1.845 ;
      RECT 6.435 0.87 6.99 1.155 ;
      RECT 4.63 1.44 4.895 1.7 ;
      RECT 4.685 1.3 4.895 1.7 ;
      RECT 4.685 0.83 4.865 1.7 ;
      RECT 3.095 0.825 3.345 1.01 ;
      RECT 3.095 0.83 4.865 0.99 ;
      RECT 3.095 0.825 3.46 0.99 ;
      RECT 1.63 3.08 2.765 3.24 ;
      RECT 2.605 2.52 2.765 3.24 ;
      RECT 3.365 2.985 4.645 3.145 ;
      RECT 4.29 2.685 4.645 3.145 ;
      RECT 1.63 2.835 1.815 3.24 ;
      RECT 0.84 2.835 1.815 2.995 ;
      RECT 3.365 2.52 3.535 3.145 ;
      RECT 0.685 0.645 0.845 2.935 ;
      RECT 0.685 2.2 1.01 2.935 ;
      RECT 4.29 1.17 4.45 3.145 ;
      RECT 2.605 2.52 3.535 2.68 ;
      RECT 3.385 1.225 3.645 1.64 ;
      RECT 3.465 1.17 4.45 1.33 ;
      RECT 0.315 0.645 0.845 0.84 ;
      RECT 2.245 2.145 2.425 2.9 ;
      RECT 3.89 1.51 4.075 2.805 ;
      RECT 2.245 2.145 4.075 2.315 ;
      RECT 1.835 2.145 4.075 2.305 ;
      RECT 1.835 1.67 2.155 2.305 ;
      RECT 3.89 1.51 4.11 1.81 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dfrbp_2

MACRO sg13g2_dlhq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlhq_1 0 0 ;
  SIZE 8.16 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.315 1.4 0.785 2.07 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.575 1.57 6.905 2 ;
    END
  END GATE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.45 2.075 7.785 3.155 ;
        RECT 7.625 0.63 7.785 3.155 ;
        RECT 7.435 0.63 7.785 1.355 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 8.16 4 ;
        RECT 6.965 2.23 7.225 4 ;
        RECT 5.03 3.115 5.305 4 ;
        RECT 1.85 3.19 2.11 4 ;
        RECT 0.275 2.4 0.535 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 8.16 0.22 ;
        RECT 6.88 -0.22 7.14 0.515 ;
        RECT 5.27 -0.22 5.55 0.445 ;
        RECT 1.925 -0.22 2.185 1.27 ;
        RECT 0.335 -0.22 0.595 1.03 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 4.5 1.93 5.005 2.195 ;
      RECT 4.77 0.475 5.005 2.195 ;
      RECT 7.085 1.54 7.445 1.87 ;
      RECT 7.085 0.7 7.255 1.87 ;
      RECT 6.29 0.7 7.255 0.88 ;
      RECT 4.77 0.625 6.5 0.785 ;
      RECT 2.39 0.475 2.665 0.78 ;
      RECT 2.39 0.475 5.005 0.635 ;
      RECT 3.78 2.725 6.715 2.885 ;
      RECT 6.035 2.205 6.715 2.885 ;
      RECT 3.78 1.93 3.95 2.885 ;
      RECT 6.035 1.57 6.395 2.885 ;
      RECT 6.235 1.115 6.395 2.885 ;
      RECT 3.39 1.93 3.95 2.095 ;
      RECT 3.045 1.655 3.545 1.975 ;
      RECT 6.235 1.115 6.6 1.39 ;
      RECT 4.13 2.385 5.815 2.545 ;
      RECT 5.565 1.005 5.815 2.545 ;
      RECT 4.13 1.515 4.29 2.545 ;
      RECT 3.735 1.515 4.29 1.75 ;
      RECT 5.565 1.005 6.055 1.265 ;
      RECT 3.05 2.275 3.6 2.435 ;
      RECT 2.705 2.155 3.205 2.315 ;
      RECT 2.705 1.315 2.865 2.315 ;
      RECT 2.705 1.315 3.545 1.475 ;
      RECT 4.255 0.995 4.585 1.325 ;
      RECT 3.225 1.155 4.585 1.325 ;
      RECT 3.33 3.065 4.175 3.235 ;
      RECT 3.33 2.615 3.5 3.235 ;
      RECT 2.71 2.615 3.5 2.785 ;
      RECT 2.27 2.495 2.865 2.66 ;
      RECT 2.27 2.225 2.52 2.66 ;
      RECT 1.535 1.575 2.525 1.745 ;
      RECT 2.365 0.965 2.525 1.745 ;
      RECT 1.535 0.725 1.695 1.745 ;
      RECT 2.365 0.965 3.02 1.13 ;
      RECT 1.415 0.725 1.695 1.035 ;
      RECT 2.85 0.815 4.02 0.975 ;
      RECT 2.355 3.025 3.04 3.205 ;
      RECT 1.335 2.215 1.57 3.165 ;
      RECT 2.355 2.84 2.525 3.205 ;
      RECT 1.335 2.84 2.525 3 ;
      RECT 0.785 2.405 1.135 3.135 ;
      RECT 0.965 1.32 1.135 3.135 ;
      RECT 0.965 1.32 1.355 1.99 ;
      RECT 0.965 0.79 1.125 3.135 ;
      RECT 0.825 0.79 1.125 1.095 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlhq_1

MACRO sg13g2_dlhr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlhr_1 0 0 ;
  SIZE 8.64 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.765 1.45 1.11 1.91 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.29 1.45 1.59 1.91 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.63 1.325 6.05 1.875 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.53 2.395 6.945 3.175 ;
        RECT 6.785 1.01 6.945 3.175 ;
        RECT 6.435 1.01 6.945 1.24 ;
        RECT 6.435 0.51 6.72 1.24 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 8.64 4 ;
        RECT 7.635 2.31 7.82 4 ;
        RECT 6.095 2.46 6.285 4 ;
        RECT 4.7 2.835 5.3 4 ;
        RECT 2.65 2.935 2.93 4 ;
        RECT 0.97 2.935 1.23 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 8.64 0.22 ;
        RECT 7.55 -0.22 7.81 1.12 ;
        RECT 5.905 -0.22 6.235 1.14 ;
        RECT 4.545 -0.22 4.83 1.115 ;
        RECT 2.645 -0.22 2.905 0.54 ;
        RECT 0.91 -0.22 1.24 1.25 ;
    END
  END VSS
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8 1.97 8.39 3.09 ;
        RECT 8.215 0.47 8.39 3.09 ;
        RECT 8.02 0.47 8.39 1.085 ;
    END
  END Q_N
  OBS
    LAYER Metal1 ;
      RECT 7.125 1.475 7.315 3.09 ;
      RECT 7.125 1.475 8 1.76 ;
      RECT 7.125 0.49 7.305 3.09 ;
      RECT 7 0.49 7.305 0.775 ;
      RECT 5.575 2.055 5.78 3.09 ;
      RECT 4.51 2.12 5.78 2.45 ;
      RECT 6.29 1.48 6.605 2.215 ;
      RECT 5.29 2.055 6.605 2.215 ;
      RECT 5.29 0.51 5.45 2.45 ;
      RECT 5.085 0.51 5.45 1.23 ;
      RECT 3.495 2.535 3.8 2.855 ;
      RECT 3.64 1.77 3.8 2.855 ;
      RECT 3.64 1.77 5.11 1.935 ;
      RECT 4.84 1.48 5.11 1.935 ;
      RECT 3.865 1.76 5.11 1.935 ;
      RECT 3.865 0.84 4.035 1.935 ;
      RECT 3.59 0.84 4.035 1.09 ;
      RECT 3.14 3.035 4.3 3.205 ;
      RECT 3.99 2.18 4.3 3.205 ;
      RECT 3.14 2.105 3.31 3.205 ;
      RECT 2.11 2.125 2.5 2.415 ;
      RECT 2.33 1.075 2.5 2.415 ;
      RECT 3.3 1.27 3.46 2.27 ;
      RECT 3.3 1.27 3.68 1.59 ;
      RECT 2.33 1.27 3.68 1.435 ;
      RECT 2.11 1.075 2.5 1.35 ;
      RECT 1.52 2.165 1.93 2.355 ;
      RECT 1.77 0.66 1.93 2.355 ;
      RECT 1.77 1.55 2.145 1.88 ;
      RECT 1.455 0.66 1.93 1.25 ;
      RECT 1.455 0.72 3.275 0.89 ;
      RECT 3.105 0.44 3.275 0.89 ;
      RECT 3.105 0.44 4.19 0.63 ;
      RECT 0.38 2.3 0.665 2.945 ;
      RECT 0.38 2.595 2.96 2.755 ;
      RECT 2.79 1.62 2.96 2.755 ;
      RECT 0.38 0.96 0.54 2.945 ;
      RECT 2.79 1.62 3.12 1.92 ;
      RECT 0.38 0.96 0.665 1.27 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlhr_1

MACRO sg13g2_dlhrq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlhrq_1 0 0 ;
  SIZE 7.2 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.52 0.6 2 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.185 1.505 1.525 2 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.695 1.57 6.015 2 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6884 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.525 2.075 6.885 3.16 ;
        RECT 6.725 0.77 6.885 3.16 ;
        RECT 6.395 0.77 6.885 1.02 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.2 4 ;
        RECT 6.025 2.205 6.23 4 ;
        RECT 4.875 2.935 5.135 4 ;
        RECT 2.62 2.935 2.88 4 ;
        RECT 0.87 2.935 1.13 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.2 0.22 ;
        RECT 5.905 -0.22 6.165 0.985 ;
        RECT 4.49 -0.22 4.75 0.895 ;
        RECT 2.59 -0.22 2.88 0.745 ;
        RECT 0.995 -0.22 1.26 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 5.495 2.205 5.735 3.16 ;
      RECT 4.555 2.3 5.735 2.585 ;
      RECT 5.355 1.2 5.515 2.585 ;
      RECT 6.225 1.2 6.545 1.77 ;
      RECT 5.025 1.2 6.545 1.36 ;
      RECT 5.025 0.64 5.285 1.36 ;
      RECT 3.545 2.66 3.785 2.92 ;
      RECT 3.625 1.945 3.785 2.92 ;
      RECT 3.625 1.955 5.175 2.115 ;
      RECT 4.915 1.69 5.175 2.115 ;
      RECT 3.745 0.85 3.905 2.115 ;
      RECT 3.535 0.85 3.905 1.085 ;
      RECT 1.465 2.18 1.875 2.415 ;
      RECT 1.705 1.68 1.875 2.415 ;
      RECT 1.705 1.68 2.08 2 ;
      RECT 4.085 1.445 4.345 1.775 ;
      RECT 1.705 0.925 1.865 2.415 ;
      RECT 4.085 0.475 4.255 1.775 ;
      RECT 1.485 0.605 1.775 1.315 ;
      RECT 1.485 0.925 3.27 1.085 ;
      RECT 3.1 0.475 3.27 1.085 ;
      RECT 3.1 0.475 4.255 0.645 ;
      RECT 3.155 3.18 4.295 3.34 ;
      RECT 3.965 2.295 4.295 3.34 ;
      RECT 3.155 2.195 3.325 3.34 ;
      RECT 2.055 2.2 2.42 2.415 ;
      RECT 2.26 1.265 2.42 2.415 ;
      RECT 3.285 1.265 3.445 2.37 ;
      RECT 3.285 1.265 3.565 1.67 ;
      RECT 2.045 1.265 3.565 1.445 ;
      RECT 0.365 2.37 0.61 3.14 ;
      RECT 0.365 2.595 2.945 2.755 ;
      RECT 2.775 1.69 2.945 2.755 ;
      RECT 0.365 2.37 0.965 2.755 ;
      RECT 0.78 1.12 0.965 2.755 ;
      RECT 2.775 1.69 3.105 2.02 ;
      RECT 0.24 1.12 0.965 1.34 ;
      RECT 0.24 0.92 0.515 1.34 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlhrq_1

MACRO sg13g2_dllr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dllr_1 0 0 ;
  SIZE 9.12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 1.48 1.1 2.12 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.29 1.49 1.61 2.12 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.11 1.41 6.45 1.81 ;
    END
  END RESET_B
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.55 2.07 8.96 3.135 ;
        RECT 8.715 0.54 8.96 3.135 ;
        RECT 8.595 0.54 8.96 1.22 ;
    END
  END Q_N
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.245 1.135 7.435 2.2 ;
        RECT 6.89 0.535 7.365 1.25 ;
        RECT 6.975 1.965 7.31 3.035 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 9.12 4 ;
        RECT 8.15 2.06 8.33 4 ;
        RECT 6.455 2.425 6.715 4 ;
        RECT 5.02 2.815 5.695 4 ;
        RECT 2.825 3.12 3.085 4 ;
        RECT 0.905 2.895 1.165 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 8.085 -0.22 9.12 0.305 ;
        RECT 8.085 -0.22 8.345 1.22 ;
        RECT 0 -0.22 9.12 0.22 ;
        RECT 6.38 -0.22 6.64 1.16 ;
        RECT 5.01 -0.22 5.24 1.165 ;
        RECT 2.785 -0.22 3.045 0.82 ;
        RECT 0.95 -0.22 1.21 1.235 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 7.53 2.355 7.825 2.96 ;
      RECT 7.615 0.725 7.825 2.96 ;
      RECT 7.615 1.52 8.52 1.85 ;
      RECT 7.615 0.725 7.835 1.85 ;
      RECT 7.545 0.725 7.835 0.98 ;
      RECT 5.9 1.99 6.23 3.07 ;
      RECT 4.815 2.2 6.23 2.51 ;
      RECT 6.635 1.48 6.795 2.245 ;
      RECT 5.605 1.99 6.795 2.245 ;
      RECT 5.605 0.555 5.78 2.51 ;
      RECT 6.635 1.48 7.06 1.77 ;
      RECT 5.495 0.555 5.78 1.27 ;
      RECT 3.785 2.625 4.075 2.955 ;
      RECT 3.915 1.855 4.075 2.955 ;
      RECT 3.915 1.855 5.01 2.02 ;
      RECT 4.67 1.44 5.01 2.02 ;
      RECT 4.67 1.44 5.405 1.77 ;
      RECT 4.67 0.595 4.83 2.02 ;
      RECT 3.835 0.595 4.83 0.83 ;
      RECT 3.405 3.155 4.55 3.34 ;
      RECT 4.275 2.27 4.55 3.34 ;
      RECT 3.405 2.2 3.575 3.34 ;
      RECT 1.69 2.43 1.96 2.695 ;
      RECT 1.69 2.43 2.84 2.59 ;
      RECT 2.67 1.35 2.84 2.59 ;
      RECT 1.69 2.41 1.95 2.695 ;
      RECT 1.79 0.595 1.95 2.695 ;
      RECT 3.565 1.35 3.735 2.365 ;
      RECT 2.505 1.465 2.84 1.77 ;
      RECT 3.565 1.35 3.895 1.67 ;
      RECT 2.52 1.35 3.895 1.51 ;
      RECT 1.51 0.595 1.95 1.29 ;
      RECT 2.13 1.955 2.485 2.25 ;
      RECT 2.13 0.605 2.3 2.25 ;
      RECT 4.16 1.01 4.49 1.67 ;
      RECT 2.13 0.605 2.38 1.225 ;
      RECT 2.13 1.01 4.49 1.17 ;
      RECT 2.13 0.605 2.39 1.17 ;
      RECT 1.35 2.95 2.3 3.12 ;
      RECT 2.13 2.78 2.3 3.12 ;
      RECT 0.38 2.355 0.655 3.12 ;
      RECT 1.35 2.355 1.51 3.12 ;
      RECT 2.13 2.78 3.195 2.94 ;
      RECT 3.025 1.69 3.195 2.94 ;
      RECT 0.38 2.355 1.51 2.515 ;
      RECT 0.38 0.875 0.54 3.12 ;
      RECT 3.025 1.69 3.355 2.02 ;
      RECT 0.38 0.875 0.66 1.185 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dllr_1

MACRO sg13g2_dllrq_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dllrq_1 0 0 ;
  SIZE 7.68 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1.56 1.115 1.96 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2054 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.305 1.56 1.62 1.96 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.13 1.29 6.535 1.915 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8449 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.085 2.085 7.415 3.155 ;
        RECT 7.255 0.5 7.415 3.155 ;
        RECT 7.065 0.5 7.415 1.2 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.68 4 ;
        RECT 6.45 2.56 6.705 4 ;
        RECT 4.975 2.7 5.655 4 ;
        RECT 2.715 3.025 2.975 4 ;
        RECT 0.99 2.155 1.25 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.68 0.22 ;
        RECT 6.475 -0.22 6.735 1.105 ;
        RECT 5.01 -0.22 5.27 0.725 ;
        RECT 2.695 -0.22 3.46 0.49 ;
        RECT 0.96 -0.22 1.22 0.49 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 5.905 2.215 6.165 3.03 ;
      RECT 5.78 0.495 5.95 2.47 ;
      RECT 4.785 2.215 6.885 2.375 ;
      RECT 6.715 1.43 6.885 2.375 ;
      RECT 4.785 2.14 5.95 2.47 ;
      RECT 6.715 1.43 7.075 1.76 ;
      RECT 5.55 0.495 5.95 1.2 ;
      RECT 3.555 2.29 4.035 2.46 ;
      RECT 3.875 1.8 4.035 2.46 ;
      RECT 3.875 1.8 5.37 1.96 ;
      RECT 5.185 1.41 5.37 1.96 ;
      RECT 5.185 1.41 5.595 1.74 ;
      RECT 5.185 0.915 5.355 1.96 ;
      RECT 4.135 0.915 5.355 1.075 ;
      RECT 4.135 0.56 4.395 1.075 ;
      RECT 2.165 2.125 2.545 2.385 ;
      RECT 2.385 1.015 2.545 2.385 ;
      RECT 2.385 1.95 3.69 2.11 ;
      RECT 3.375 1.3 3.69 2.11 ;
      RECT 3.375 1.3 4.635 1.615 ;
      RECT 2.145 1.015 2.545 1.28 ;
      RECT 1.49 2.68 1.975 2.855 ;
      RECT 1.49 2.68 4.545 2.84 ;
      RECT 4.215 2.14 4.545 2.84 ;
      RECT 1.49 2.14 1.965 2.855 ;
      RECT 1.805 1.07 1.965 2.855 ;
      RECT 1.805 1.46 2.205 1.78 ;
      RECT 1.495 1.07 1.965 1.335 ;
      RECT 0.395 2.14 0.75 2.855 ;
      RECT 0.395 0.67 0.565 2.855 ;
      RECT 2.835 0.67 3.165 1.7 ;
      RECT 0.395 0.67 0.745 1.36 ;
      RECT 0.395 0.67 3.165 0.835 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dllrq_1

MACRO sg13g2_dlygate4sd1_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlygate4sd1_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.425 0.835 1.945 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.43 2.075 3.72 3.16 ;
        RECT 3.455 0.61 3.72 3.16 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.9 2.455 3.16 4 ;
        RECT 0.745 2.665 1.01 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.915 -0.22 3.175 0.965 ;
        RECT 0.69 -0.22 1.02 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.14 2.03 2.45 2.395 ;
      RECT 2.14 2.03 3.235 2.205 ;
      RECT 3.045 1.16 3.235 2.205 ;
      RECT 3.045 1.16 3.265 1.845 ;
      RECT 2.155 1.16 3.265 1.36 ;
      RECT 2.155 0.96 2.395 1.36 ;
      RECT 1.52 2.615 1.825 2.945 ;
      RECT 1.58 1.57 1.825 2.945 ;
      RECT 1.58 1.57 2.79 1.83 ;
      RECT 1.58 0.665 1.81 2.945 ;
      RECT 1.52 0.665 1.81 0.95 ;
      RECT 0.24 2.195 0.5 2.91 ;
      RECT 0.24 2.195 1.375 2.4 ;
      RECT 1.12 1.065 1.375 2.4 ;
      RECT 0.21 1.065 1.375 1.24 ;
      RECT 0.21 0.66 0.48 1.24 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlygate4sd1_1

MACRO sg13g2_dlygate4sd2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlygate4sd2_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.425 0.835 1.945 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.43 2.075 3.72 3.16 ;
        RECT 3.455 0.61 3.72 3.16 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.9 2.455 3.16 4 ;
        RECT 0.745 2.665 1.01 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.915 -0.22 3.175 0.965 ;
        RECT 0.69 -0.22 1.02 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.14 2.03 2.45 2.395 ;
      RECT 2.14 2.03 3.235 2.205 ;
      RECT 3.045 1.16 3.235 2.205 ;
      RECT 3.045 1.16 3.265 1.845 ;
      RECT 2.155 1.16 3.265 1.36 ;
      RECT 2.155 0.96 2.395 1.36 ;
      RECT 1.52 2.615 1.825 2.945 ;
      RECT 1.58 1.57 1.825 2.945 ;
      RECT 1.58 1.57 2.79 1.83 ;
      RECT 1.58 0.665 1.81 2.945 ;
      RECT 1.52 0.665 1.81 0.95 ;
      RECT 0.24 2.195 0.5 2.91 ;
      RECT 0.24 2.195 1.375 2.4 ;
      RECT 1.12 1.065 1.375 2.4 ;
      RECT 0.21 1.065 1.375 1.24 ;
      RECT 0.21 0.66 0.48 1.24 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlygate4sd2_1

MACRO sg13g2_dlygate4sd3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_dlygate4sd3_1 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1092 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 1.41 0.915 2.08 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 3.1 2.395 3.36 4 ;
        RECT 0.81 2.665 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 3.13 -0.22 3.39 0.85 ;
        RECT 0.8 -0.22 1.07 0.835 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 2.075 4.02 3.17 ;
        RECT 3.805 0.595 4.02 3.17 ;
        RECT 3.61 0.595 4.02 1.34 ;
    END
  END X
  OBS
    LAYER Metal1 ;
      RECT 2.205 2.045 2.465 2.38 ;
      RECT 2.205 2.045 3.34 2.215 ;
      RECT 3.15 1.045 3.34 2.215 ;
      RECT 3.15 1.515 3.535 1.845 ;
      RECT 2.205 1.045 3.34 1.235 ;
      RECT 2.205 0.945 2.47 1.235 ;
      RECT 1.675 2.615 1.955 2.93 ;
      RECT 1.72 0.665 1.955 2.93 ;
      RECT 1.72 1.55 2.925 1.81 ;
      RECT 0.3 2.32 0.56 2.88 ;
      RECT 0.3 2.32 1.455 2.48 ;
      RECT 1.175 1.015 1.455 2.48 ;
      RECT 0.3 1.015 1.455 1.205 ;
      RECT 0.3 0.69 0.56 1.205 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_dlygate4sd3_1

MACRO sg13g2_ebufn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_ebufn_2 0 0 ;
  SIZE 4.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.5044 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 1.37 3.495 1.85 ;
    END
  END TE_B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.695 1.52 4.055 1.925 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.94 1.965 2.26 ;
        RECT 0.84 1.94 1.1 2.61 ;
        RECT 0.74 0.845 1.025 1.08 ;
        RECT 0.74 0.845 0.91 2.14 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.8 4 ;
        RECT 3.52 2.895 3.78 4 ;
        RECT 1.89 3.18 2.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.8 0.22 ;
        RECT 3.56 -0.22 3.82 1.13 ;
        RECT 1.78 -0.22 2.04 0.88 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 4.14 2.085 4.435 2.95 ;
      RECT 4.245 0.595 4.435 2.95 ;
      RECT 2.155 2.495 4.435 2.66 ;
      RECT 2.155 1.485 2.325 2.66 ;
      RECT 1.09 1.485 2.325 1.75 ;
      RECT 4.06 0.595 4.435 1.13 ;
      RECT 2.7 2.035 3.295 2.3 ;
      RECT 2.7 0.525 2.915 2.3 ;
      RECT 2.7 0.525 3.3 1.18 ;
      RECT 0.33 3.075 1.61 3.32 ;
      RECT 1.35 2.52 1.61 3.32 ;
      RECT 2.435 2.84 2.705 3.13 ;
      RECT 0.33 2.395 0.59 3.32 ;
      RECT 1.35 2.84 2.705 3 ;
      RECT 1.28 1.13 2.515 1.3 ;
      RECT 2.3 0.54 2.515 1.3 ;
      RECT 0.25 0.44 0.51 1.215 ;
      RECT 1.28 0.44 1.505 1.3 ;
      RECT 0.25 0.44 1.505 0.635 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_ebufn_2

MACRO sg13g2_ebufn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_ebufn_4 0 0 ;
  SIZE 6.72 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.5 0.99 1.95 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8242 LAYER Metal1 ;
      ANTENNAGATEAREA 0.8242 LAYER Metal2 ;
      ANTENNAMAXAREACAR 0.152633 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.0438 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.17 1.33 1.51 1.7 ;
      LAYER Metal2 ;
        RECT 1.3 1.345 1.59 1.95 ;
      LAYER Via1 ;
        RECT 1.305 1.435 1.495 1.625 ;
    END
  END TE_B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4322 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.75 2.11 6.01 2.765 ;
        RECT 5.83 0.95 6.01 2.765 ;
        RECT 4.715 1.145 6.01 1.375 ;
        RECT 5.745 0.95 6.01 1.375 ;
        RECT 4.72 2.11 6.01 2.335 ;
        RECT 4.72 2.11 4.98 2.885 ;
        RECT 4.715 0.95 4.975 1.375 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 6.72 4 ;
        RECT 3.69 2.455 3.95 4 ;
        RECT 2.67 2.945 2.93 4 ;
        RECT 0.89 2.915 1.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 6.72 0.22 ;
        RECT 3.69 -0.22 3.95 0.895 ;
        RECT 2.67 -0.22 2.93 1.145 ;
        RECT 0.805 -0.22 1.065 1.15 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.19 1.325 3.44 1.485 ;
      RECT 3.18 0.62 3.44 1.485 ;
      RECT 4.24 0.455 4.42 1.425 ;
      RECT 3.18 1.23 4.42 1.425 ;
      RECT 2.19 0.57 2.385 1.485 ;
      RECT 6.26 0.455 6.52 1.245 ;
      RECT 5.235 0.455 5.495 0.88 ;
      RECT 4.24 0.455 6.52 0.625 ;
      RECT 4.245 3.17 6.52 3.33 ;
      RECT 6.26 2.165 6.52 3.33 ;
      RECT 5.24 2.585 5.5 3.33 ;
      RECT 4.245 2.115 4.415 3.33 ;
      RECT 3.18 2.115 3.44 3.13 ;
      RECT 2.19 2.6 2.46 3.05 ;
      RECT 2.19 2.6 3.44 2.765 ;
      RECT 3.18 2.115 4.415 2.275 ;
      RECT 0.28 2.15 0.635 3.17 ;
      RECT 0.28 2.57 2.01 2.73 ;
      RECT 1.815 2.26 2.01 2.73 ;
      RECT 2.63 1.7 2.8 2.39 ;
      RECT 1.87 2.23 2.8 2.39 ;
      RECT 0.28 0.59 0.445 3.17 ;
      RECT 2.63 1.7 5.57 1.86 ;
      RECT 4.575 1.555 5.57 1.86 ;
      RECT 0.28 0.59 0.525 1.31 ;
      RECT 1.41 1.9 1.635 2.39 ;
      RECT 1.41 1.9 1.755 2.09 ;
      RECT 1.75 0.5 2.01 2.04 ;
      RECT 1.58 1.87 2.01 2.04 ;
      RECT 1.315 0.5 2.01 1.15 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_ebufn_4

MACRO sg13g2_ebufn_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_ebufn_8 0 0 ;
  SIZE 12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8272 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.73 2.12 3.99 2.85 ;
        RECT 0.67 1.17 3.99 1.36 ;
        RECT 3.73 0.915 3.99 1.36 ;
        RECT 0.67 2.12 3.99 2.29 ;
        RECT 2.71 2.12 2.97 2.86 ;
        RECT 2.71 0.92 2.97 1.36 ;
        RECT 0.67 2.12 2.97 2.295 ;
        RECT 1.69 2.12 1.95 2.83 ;
        RECT 1.685 0.92 1.95 1.36 ;
        RECT 0.78 1.17 1.14 2.295 ;
        RECT 0.67 2.02 0.93 2.82 ;
        RECT 0.67 0.92 0.93 1.465 ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.84 1.455 11.335 1.835 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.4066 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.61 1.51 10.63 1.835 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 12 4 ;
        RECT 11.51 2.62 11.77 4 ;
        RECT 10.49 2.915 10.75 4 ;
        RECT 7.84 3.205 8.105 4 ;
        RECT 6.795 2.975 7.055 4 ;
        RECT 5.77 2.96 6.03 4 ;
        RECT 4.75 2.97 5.01 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 12 0.22 ;
        RECT 11.51 -0.22 11.77 0.855 ;
        RECT 10.49 -0.22 10.75 1.22 ;
        RECT 7.875 -0.22 8.135 1.225 ;
        RECT 6.855 -0.22 7.115 1.225 ;
        RECT 5.835 -0.22 6.095 1.225 ;
        RECT 4.815 -0.22 5.075 1.2 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 11 2.24 11.26 3.155 ;
      RECT 8.805 2.56 11.26 2.725 ;
      RECT 8.805 2.25 8.985 2.725 ;
      RECT 11 2.24 11.765 2.44 ;
      RECT 11.59 1.09 11.765 2.44 ;
      RECT 4.235 2.25 8.985 2.41 ;
      RECT 4.235 1.73 4.445 2.41 ;
      RECT 1.58 1.73 4.445 1.9 ;
      RECT 1.58 1.585 3.995 1.9 ;
      RECT 11 1.09 11.765 1.26 ;
      RECT 11 0.675 11.26 1.26 ;
      RECT 9.165 2.1 10.24 2.38 ;
      RECT 9.165 0.59 9.4 2.38 ;
      RECT 9.165 0.59 10.24 1.22 ;
      RECT 8.855 0.59 10.24 0.92 ;
      RECT 0.16 3.155 4.495 3.325 ;
      RECT 4.27 2.59 4.495 3.325 ;
      RECT 8.365 2.84 8.665 3.23 ;
      RECT 7.305 2.59 7.565 3.16 ;
      RECT 6.285 2.59 6.55 3.16 ;
      RECT 5.26 2.59 5.52 3.155 ;
      RECT 3.22 2.47 3.48 3.325 ;
      RECT 2.2 2.48 2.46 3.325 ;
      RECT 1.18 2.48 1.44 3.325 ;
      RECT 0.16 2.15 0.42 3.325 ;
      RECT 7.305 2.84 8.665 3.02 ;
      RECT 6.285 2.59 7.565 2.79 ;
      RECT 4.27 2.59 7.565 2.78 ;
      RECT 4.72 1.55 8.645 1.72 ;
      RECT 8.385 0.675 8.645 1.72 ;
      RECT 4.28 1.38 5.585 1.55 ;
      RECT 7.365 0.68 7.625 1.72 ;
      RECT 6.345 0.675 6.605 1.72 ;
      RECT 5.325 0.68 5.585 1.72 ;
      RECT 4.28 0.53 4.525 1.55 ;
      RECT 0.15 0.53 0.405 1.34 ;
      RECT 3.22 0.53 3.48 0.985 ;
      RECT 2.2 0.53 2.46 0.985 ;
      RECT 1.18 0.53 1.44 0.975 ;
      RECT 0.15 0.53 4.525 0.73 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_ebufn_8

MACRO sg13g2_einvn_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_einvn_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.16 1.005 3.49 2.945 ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.7 1.01 4.03 1.75 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.429 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.28 1.32 0.995 2.33 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 2.14 2.43 2.4 4 ;
        RECT 0.6 2.745 0.86 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 2.15 -0.22 2.41 0.915 ;
        RECT 0.625 -0.22 0.875 0.96 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.655 1.095 2.92 1.305 ;
      RECT 2.665 0.55 2.92 1.305 ;
      RECT 1.655 0.575 1.9 1.305 ;
      RECT 2.665 0.55 3.95 0.825 ;
      RECT 2.685 3.175 3.93 3.335 ;
      RECT 3.67 2.11 3.93 3.335 ;
      RECT 2.685 2.045 2.875 3.335 ;
      RECT 1.645 2.045 1.895 3.145 ;
      RECT 1.645 2.045 2.875 2.235 ;
      RECT 1.085 2.745 1.385 3.14 ;
      RECT 1.215 0.595 1.385 3.14 ;
      RECT 1.215 1.52 1.655 1.85 ;
      RECT 1.085 0.595 1.385 0.96 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_einvn_2

MACRO sg13g2_einvn_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_einvn_4 0 0 ;
  SIZE 6.24 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.2 1.025 5.565 1.205 ;
        RECT 5.295 0.915 5.565 1.205 ;
        RECT 5.1 2.13 5.36 2.955 ;
        RECT 4.08 2.13 5.36 2.33 ;
        RECT 4.2 1.025 4.435 2.33 ;
        RECT 4.08 2.015 4.34 2.955 ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9672 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.615 1.44 5.735 1.91 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8242 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.46 0.695 2 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 6.24 4 ;
        RECT 3.06 2.245 3.32 4 ;
        RECT 2.04 2.25 2.3 4 ;
        RECT 0.365 2.21 0.625 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 6.24 0.22 ;
        RECT 3.26 -0.22 3.52 1.185 ;
        RECT 2.24 -0.22 2.5 1.195 ;
        RECT 0.4 -0.22 0.67 1.205 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.77 1.385 4 1.575 ;
      RECT 3.8 0.605 4 1.575 ;
      RECT 2.75 0.74 3.01 1.575 ;
      RECT 1.77 0.57 1.965 1.575 ;
      RECT 5.81 0.475 6.07 0.99 ;
      RECT 3.8 0.605 5.06 0.84 ;
      RECT 4.77 0.475 6.07 0.645 ;
      RECT 3.61 3.14 5.87 3.335 ;
      RECT 5.61 2.115 5.87 3.335 ;
      RECT 4.59 2.54 4.85 3.335 ;
      RECT 3.61 1.795 3.79 3.335 ;
      RECT 1.53 1.795 1.79 3.13 ;
      RECT 2.55 1.795 2.81 3.005 ;
      RECT 1.53 1.795 3.79 2.01 ;
      RECT 0.875 0.52 1.135 3.13 ;
      RECT 0.875 0.52 1.57 1.53 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_einvn_4

MACRO sg13g2_einvn_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_einvn_8 0 0 ;
  SIZE 10.56 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.9344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.43 1.51 9.84 1.845 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8272 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.33 2.12 9.59 2.815 ;
        RECT 6.26 1.09 9.59 1.28 ;
        RECT 9.33 0.915 9.59 1.28 ;
        RECT 6.26 2.12 9.59 2.31 ;
        RECT 8.31 2.12 8.57 2.815 ;
        RECT 8.31 0.925 8.57 1.28 ;
        RECT 7.29 2.12 7.55 2.815 ;
        RECT 7.29 1.055 7.55 1.28 ;
        RECT 6.26 1.09 6.955 2.31 ;
        RECT 6.26 1.055 6.525 2.77 ;
    END
  END Z
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.4066 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.37 0.63 1.82 ;
    END
  END TE_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 10.56 4 ;
        RECT 4.985 2.565 5.245 4 ;
        RECT 3.965 2.245 4.225 4 ;
        RECT 2.945 2.245 3.205 4 ;
        RECT 1.925 2.245 2.185 4 ;
        RECT 0.35 2.08 0.61 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 10.56 0.22 ;
        RECT 5.25 -0.22 5.51 1.21 ;
        RECT 4.23 -0.22 4.49 1.3 ;
        RECT 3.21 -0.22 3.47 1.3 ;
        RECT 2.19 -0.22 2.45 1.3 ;
        RECT 0.355 -0.22 0.615 1.18 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.72 1.49 6.005 1.66 ;
      RECT 5.765 0.57 6.005 1.66 ;
      RECT 4.74 0.665 5 1.66 ;
      RECT 3.72 0.67 3.98 1.66 ;
      RECT 2.7 0.67 2.96 1.66 ;
      RECT 1.72 0.615 1.93 1.66 ;
      RECT 9.84 0.445 10.1 1.305 ;
      RECT 8.82 0.445 9.08 0.9 ;
      RECT 7.8 0.445 8.06 0.885 ;
      RECT 6.78 0.57 7.04 0.855 ;
      RECT 5.765 0.57 8.06 0.79 ;
      RECT 7.795 0.445 10.1 0.615 ;
      RECT 5.75 3.085 10.1 3.295 ;
      RECT 9.84 2.245 10.1 3.295 ;
      RECT 1.41 1.885 1.67 3.13 ;
      RECT 4.475 2.17 4.735 3.12 ;
      RECT 3.455 1.885 3.715 3.12 ;
      RECT 2.435 1.885 2.695 3.12 ;
      RECT 8.82 2.575 9.08 3.295 ;
      RECT 7.8 2.55 8.06 3.295 ;
      RECT 6.78 2.58 7.045 3.295 ;
      RECT 5.75 2.17 6.025 3.295 ;
      RECT 4.475 2.17 6.025 2.34 ;
      RECT 4.475 1.885 4.69 3.12 ;
      RECT 1.41 1.885 4.69 2.055 ;
      RECT 0.86 1.32 1.12 3.13 ;
      RECT 0.88 0.575 1.52 1.525 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_einvn_8

MACRO sg13g2_fill_1
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_1 0 0 ;
  SIZE 0.48 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 0.48 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 0.48 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_1

MACRO sg13g2_fill_2
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_2 0 0 ;
  SIZE 0.96 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 0.96 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 0.96 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_2

MACRO sg13g2_fill_4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_4 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_4

MACRO sg13g2_fill_8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_fill_8 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_fill_8

MACRO sg13g2_inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_1 0 0 ;
  SIZE 1.44 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.44 4 ;
        RECT 0.505 2.205 0.78 4 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.651 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.045 0.595 1.275 3.175 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 1.52 0.815 2 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.44 0.22 ;
        RECT 0.485 -0.22 0.785 1.295 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_1

MACRO sg13g2_inv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_16 0 0 ;
  SIZE 9.12 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 3.8688 LAYER Metal1 ;
      ANTENNAGATEAREA 3.8688 LAYER Metal2 ;
      ANTENNAMAXAREACAR 0.036807 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.009331 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.445 1.455 7.765 1.9 ;
        RECT 6.405 1.455 6.74 1.9 ;
        RECT 5.395 1.455 5.71 1.9 ;
        RECT 4.4 1.455 4.68 1.9 ;
        RECT 3.38 1.455 3.655 1.9 ;
        RECT 2.35 1.455 2.64 1.9 ;
        RECT 1.31 1.455 1.62 1.9 ;
      LAYER Metal2 ;
        RECT 1.31 1.58 7.865 1.78 ;
      LAYER Via1 ;
        RECT 1.37 1.585 1.56 1.775 ;
        RECT 2.4 1.585 2.59 1.775 ;
        RECT 3.42 1.585 3.61 1.775 ;
        RECT 4.44 1.585 4.63 1.775 ;
        RECT 5.46 1.585 5.65 1.775 ;
        RECT 6.48 1.585 6.67 1.775 ;
        RECT 7.5 1.585 7.69 1.775 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNADIFFAREA 0.7068 LAYER Metal1 ;
    ANTENNADIFFAREA 5.6544 LAYER Metal2 ;
    PORT
      LAYER Metal1 ;
        RECT 7.975 0.625 8.235 3.14 ;
        RECT 6.955 0.625 7.215 3.14 ;
        RECT 5.935 0.625 6.195 3.135 ;
        RECT 4.915 0.625 5.175 3.13 ;
        RECT 3.895 0.625 4.155 3.13 ;
        RECT 2.875 0.625 3.135 3.125 ;
        RECT 1.855 0.63 2.115 3.125 ;
        RECT 0.835 0.63 1.095 3.135 ;
      LAYER Metal2 ;
        RECT 0.815 2 8.25 2.2 ;
      LAYER Via1 ;
        RECT 0.87 2.005 1.06 2.195 ;
        RECT 1.89 2.005 2.08 2.195 ;
        RECT 2.915 2.005 3.105 2.195 ;
        RECT 3.93 2.005 4.12 2.195 ;
        RECT 4.95 2.005 5.14 2.195 ;
        RECT 5.97 2.005 6.16 2.195 ;
        RECT 6.99 2.005 7.18 2.195 ;
        RECT 8.01 2.005 8.2 2.195 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 9.12 4 ;
        RECT 7.465 3.555 8.745 4 ;
        RECT 8.485 2.11 8.745 4 ;
        RECT 7.465 2.22 7.725 4 ;
        RECT 6.445 2.22 6.705 4 ;
        RECT 5.425 2.23 5.685 4 ;
        RECT 4.405 2.22 4.665 4 ;
        RECT 3.385 2.225 3.645 4 ;
        RECT 2.365 2.21 2.625 4 ;
        RECT 1.345 2.205 1.605 4 ;
        RECT 0.325 2.105 0.585 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 9.12 0.22 ;
        RECT 8.485 -0.22 8.745 1.27 ;
        RECT 7.465 -0.22 7.725 1.27 ;
        RECT 6.445 -0.22 6.705 1.27 ;
        RECT 5.425 -0.22 5.685 1.27 ;
        RECT 4.405 -0.22 4.665 1.27 ;
        RECT 3.385 -0.22 3.645 1.27 ;
        RECT 2.365 -0.22 2.625 1.275 ;
        RECT 1.345 -0.22 1.605 1.275 ;
        RECT 0.325 -0.22 0.585 1.28 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_16

MACRO sg13g2_inv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_2 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7124 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 0.57 1.02 3.18 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.18 1.52 0.635 2 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 1.32 2.095 1.535 4 ;
        RECT 0.275 2.185 0.535 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 1.34 -0.22 1.54 1.305 ;
        RECT 0.285 -0.22 0.545 1.3 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_2

MACRO sg13g2_inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_4 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9672 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 1.57 2 1.95 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 2.17 2.475 2.34 ;
        RECT 2.245 1.145 2.475 2.34 ;
        RECT 0.815 1.145 2.475 1.34 ;
        RECT 1.805 0.595 2.06 1.34 ;
        RECT 1.815 2.17 2.03 3.175 ;
        RECT 0.8 2.17 1.015 3.18 ;
        RECT 0.815 0.57 1.01 1.34 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.32 2.54 2.55 4 ;
        RECT 1.3 2.53 1.54 4 ;
        RECT 0.285 2.19 0.53 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.21 2.88 0.21 ;
        RECT 2.305 -0.21 2.565 0.95 ;
        RECT 1.28 -0.21 2.565 0.22 ;
        RECT 1.28 -0.21 1.55 0.945 ;
        RECT 0.27 -0.21 0.52 1.325 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_4

MACRO sg13g2_inv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_inv_8 0 0 ;
  SIZE 4.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.8458 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.74 1.42 4.44 1.84 ;
        RECT 3.775 0.64 4.035 3.19 ;
        RECT 2.74 1.18 3.015 3.2 ;
        RECT 2.755 0.665 3.015 3.2 ;
        RECT 0.715 2.22 3.015 2.38 ;
        RECT 0.715 1.18 3.015 1.345 ;
        RECT 1.735 0.635 2 1.345 ;
        RECT 1.73 2.22 1.995 3.155 ;
        RECT 0.715 2.22 1.995 2.385 ;
        RECT 0.715 2.22 0.98 3.16 ;
        RECT 0.715 0.62 0.98 1.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.9344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 1.57 2.495 2 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.8 4 ;
        RECT 4.32 2.065 4.53 4 ;
        RECT 3.29 2.055 3.5 4 ;
        RECT 2.245 2.56 2.515 4 ;
        RECT 1.215 2.565 1.495 4 ;
        RECT 0.24 2.06 0.435 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.8 0.22 ;
        RECT 4.295 -0.22 4.555 1.225 ;
        RECT 3.265 -0.22 3.525 1.195 ;
        RECT 2.245 -0.22 2.505 0.99 ;
        RECT 1.225 -0.22 1.485 1 ;
        RECT 0.205 -0.22 0.465 1.27 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_inv_8

MACRO sg13g2_lgcp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_lgcp_1 0 0 ;
  SIZE 7.2 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 1.68 1.635 2.21 ;
    END
  END GATE
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3978 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.685 1.685 5.395 2.015 ;
        RECT 5.195 1.575 5.395 2.015 ;
        RECT 4.685 1.685 4.885 2.42 ;
    END
  END CLK
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.495 1.76 6.845 3.2 ;
        RECT 6.59 0.56 6.845 3.2 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 7.2 4 ;
        RECT 5.99 2.2 6.25 4 ;
        RECT 4.72 2.73 4.98 4 ;
        RECT 3.115 3.095 3.38 4 ;
        RECT 0.89 2.89 1.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 7.2 0.22 ;
        RECT 6.09 -0.22 6.35 1.26 ;
        RECT 4.69 -0.22 4.95 1.445 ;
        RECT 2.99 0.895 3.525 1.125 ;
        RECT 3.365 -0.22 3.525 1.125 ;
        RECT 0.9 -0.22 1.115 0.8 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 5.23 2.195 5.49 2.97 ;
      RECT 5.23 2.195 5.765 2.355 ;
      RECT 5.585 0.815 5.765 2.355 ;
      RECT 5.585 1.51 6.275 1.84 ;
      RECT 5.585 0.815 5.855 1.84 ;
      RECT 5.525 0.815 5.855 1.41 ;
      RECT 4.205 2.155 4.47 2.975 ;
      RECT 3.115 2.695 4.47 2.905 ;
      RECT 3.115 1.725 3.29 2.905 ;
      RECT 1.975 2.305 3.29 2.565 ;
      RECT 1.975 1.36 2.235 2.565 ;
      RECT 4.205 1.23 4.445 2.975 ;
      RECT 3.115 1.725 3.655 2.04 ;
      RECT 3.65 2.26 4.015 2.45 ;
      RECT 3.845 0.845 4.015 2.45 ;
      RECT 2.445 1.37 2.775 2.05 ;
      RECT 2.445 1.37 4.015 1.54 ;
      RECT 3.705 0.845 4.015 1.54 ;
      RECT 0.335 2.125 0.65 3.11 ;
      RECT 0.335 0.6 0.495 3.11 ;
      RECT 0.335 0.6 0.595 1.3 ;
      RECT 0.335 0.98 1.455 1.16 ;
      RECT 1.295 0.465 1.455 1.16 ;
      RECT 2.865 0.465 3.185 0.71 ;
      RECT 1.295 0.465 3.185 0.635 ;
      RECT 1.625 2.795 2.35 3.055 ;
      RECT 1.625 2.42 1.785 3.055 ;
      RECT 0.855 2.42 1.785 2.58 ;
      RECT 0.855 1.34 1.025 2.58 ;
      RECT 0.675 1.51 1.025 1.84 ;
      RECT 0.855 1.34 1.795 1.5 ;
      RECT 1.635 0.89 1.795 1.5 ;
      RECT 1.635 0.89 2.395 1.14 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_lgcp_1

MACRO sg13g2_mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_mux2_1 0 0 ;
  SIZE 4.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.09 1.4 2.48 1.785 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.695 1.03 2.99 1.785 ;
        RECT 1.71 1.03 2.99 1.2 ;
        RECT 1.61 1.44 1.89 1.755 ;
        RECT 1.71 1.03 1.89 1.755 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 1.5 1.09 1.905 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0081 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.135 2.04 4.685 3.2 ;
        RECT 4.515 0.57 4.685 3.2 ;
        RECT 4.315 0.57 4.685 1.315 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.8 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.64 1.235 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.8 0.22 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.31 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.3 1.965 2.56 2.875 ;
      RECT 1.82 1.965 2.56 2.145 ;
      RECT 1.27 1.955 1.89 2.12 ;
      RECT 1.27 0.61 1.43 2.12 ;
      RECT 3.945 1.52 4.245 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.27 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.3 1.64 3.295 ;
      RECT 0.145 2.17 0.575 2.845 ;
      RECT 0.145 2.3 1.64 2.46 ;
      RECT 0.145 0.92 0.35 2.845 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.145 0.92 0.575 1.18 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_mux2_1

MACRO sg13g2_mux2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_mux2_2 0 0 ;
  SIZE 5.28 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.09 1.4 2.48 1.785 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2262 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.695 1.03 2.99 1.785 ;
        RECT 1.71 1.03 2.99 1.2 ;
        RECT 1.61 1.44 1.89 1.755 ;
        RECT 1.71 1.03 1.89 1.755 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 1.5 1.09 1.905 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.023 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.135 2.04 4.685 3.2 ;
        RECT 4.515 0.57 4.685 3.2 ;
        RECT 4.315 0.57 4.685 1.315 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 5.28 4 ;
        RECT 4.905 2.08 5.105 4 ;
        RECT 3.63 2.08 3.83 4 ;
        RECT 0.975 2.64 1.235 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 5.28 0.22 ;
        RECT 4.875 -0.22 5.135 1.31 ;
        RECT 3.6 -0.22 3.86 0.845 ;
        RECT 0.855 -0.22 1.09 1.31 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.3 1.965 2.56 2.875 ;
      RECT 1.825 1.965 2.56 2.135 ;
      RECT 1.27 1.95 1.91 2.12 ;
      RECT 1.27 0.61 1.43 2.12 ;
      RECT 3.945 1.52 4.245 1.85 ;
      RECT 3.945 1.03 4.135 1.85 ;
      RECT 3.195 1.03 4.135 1.2 ;
      RECT 3.195 0.61 3.365 1.2 ;
      RECT 1.27 0.61 3.365 0.83 ;
      RECT 1.48 3.125 3.425 3.295 ;
      RECT 3.25 1.54 3.425 3.295 ;
      RECT 1.48 2.3 1.64 3.295 ;
      RECT 0.145 2.17 0.575 2.845 ;
      RECT 0.145 2.3 1.64 2.46 ;
      RECT 0.145 0.92 0.35 2.845 ;
      RECT 3.25 1.54 3.72 1.87 ;
      RECT 0.145 0.92 0.575 1.18 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_mux2_2

MACRO sg13g2_mux4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_mux4_1 0 0 ;
  SIZE 10.08 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6396 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.435 1.04 1.92 ;
    END
  END S0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 1.435 1.57 1.92 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.22 1.435 3.54 2.37 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.72 1.435 4.09 2.37 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.07 1.56 6.4 2 ;
    END
  END A3
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4264 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.535 1.565 8.955 1.985 ;
    END
  END S1
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.64 2.78 9.905 3.075 ;
        RECT 9.665 0.62 9.905 3.075 ;
        RECT 9.475 0.62 9.905 1.36 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 10.08 4 ;
        RECT 9.095 2.585 9.355 4 ;
        RECT 5.95 2.905 6.28 4 ;
        RECT 3.52 2.97 3.78 4 ;
        RECT 0.985 2.12 1.245 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 10.08 0.22 ;
        RECT 9.035 -0.22 9.295 1.325 ;
        RECT 5.545 -0.22 5.805 1.01 ;
        RECT 3.495 -0.22 3.77 0.835 ;
        RECT 0.985 -0.22 1.245 0.84 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 7.01 3.125 8.91 3.295 ;
      RECT 8.75 2.23 8.91 3.295 ;
      RECT 7.01 1.335 7.3 3.295 ;
      RECT 8.75 2.23 9.46 2.4 ;
      RECT 9.195 1.57 9.46 2.4 ;
      RECT 6.965 1.16 7.21 1.505 ;
      RECT 8.195 2.17 8.57 2.92 ;
      RECT 8.195 0.755 8.355 2.92 ;
      RECT 7.85 1.665 8.355 1.995 ;
      RECT 8.195 0.755 8.745 1.385 ;
      RECT 4.525 2.2 5.385 2.945 ;
      RECT 7.51 2.22 7.86 2.92 ;
      RECT 4.525 2.2 5.885 2.37 ;
      RECT 5.715 1.21 5.885 2.37 ;
      RECT 7.51 1.325 7.67 2.92 ;
      RECT 7.51 1.325 8.015 1.485 ;
      RECT 7.855 0.44 8.015 1.485 ;
      RECT 5.15 1.21 6.375 1.38 ;
      RECT 6.115 0.44 6.375 1.38 ;
      RECT 5.15 0.595 5.32 1.38 ;
      RECT 4.55 0.595 5.32 0.87 ;
      RECT 6.115 0.44 8.015 0.6 ;
      RECT 4.015 3.125 5.77 3.295 ;
      RECT 5.57 2.555 5.77 3.295 ;
      RECT 6.51 2.17 6.78 3.2 ;
      RECT 6.58 0.82 6.78 3.2 ;
      RECT 4.015 2.555 4.24 3.295 ;
      RECT 2.26 1.95 2.77 2.905 ;
      RECT 5.57 2.555 6.78 2.725 ;
      RECT 2.26 2.555 4.24 2.725 ;
      RECT 2.26 0.87 2.42 2.905 ;
      RECT 2.095 0.87 2.42 1.2 ;
      RECT 7.45 0.82 7.675 1.08 ;
      RECT 6.58 0.82 7.675 0.98 ;
      RECT 0.33 2.12 0.745 2.985 ;
      RECT 0.33 0.59 0.5 2.985 ;
      RECT 4.8 1.665 5.535 1.97 ;
      RECT 1.75 1.42 2.08 1.75 ;
      RECT 4.3 1.05 4.61 1.67 ;
      RECT 2.68 1.05 3.01 1.67 ;
      RECT 4.8 1.05 4.97 1.97 ;
      RECT 1.75 0.475 1.915 1.75 ;
      RECT 2.68 1.05 4.97 1.21 ;
      RECT 0.33 1.02 1.915 1.2 ;
      RECT 2.68 0.475 2.85 1.67 ;
      RECT 0.33 0.59 0.64 1.2 ;
      RECT 1.75 0.475 2.85 0.645 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_mux4_1

MACRO sg13g2_nand2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2_1 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 1.06 1.475 1.245 ;
        RECT 1.215 0.655 1.475 1.245 ;
        RECT 0.83 1.365 1.09 3.125 ;
        RECT 0.86 1.06 1.09 3.125 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.27 1.44 1.6 1.81 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 1.44 0.62 1.81 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 1.34 2.125 1.6 4 ;
        RECT 0.32 2.125 0.58 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.395 -0.22 0.655 1.245 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2_1

MACRO sg13g2_nand2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1248 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 2.16 2.15 3.18 ;
        RECT 1.38 1.39 2.14 1.55 ;
        RECT 1.88 1 2.14 1.55 ;
        RECT 0.84 2.16 2.15 2.36 ;
        RECT 0.84 2.14 1.62 2.36 ;
        RECT 1.38 1.39 1.62 2.36 ;
        RECT 0.84 2.14 1.1 3.18 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.73 2.645 1.98 ;
        RECT 2.37 1.44 2.645 1.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 1.39 1.15 1.92 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.39 2.16 2.65 4 ;
        RECT 1.35 2.9 1.61 4 ;
        RECT 0.32 2.125 0.58 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 0.85 -0.22 1.11 0.855 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.37 0.53 2.65 1.2 ;
      RECT 0.325 1.035 1.62 1.2 ;
      RECT 1.35 0.53 1.62 1.2 ;
      RECT 0.325 0.5 0.585 1.2 ;
      RECT 1.35 0.53 2.65 0.76 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2_2

MACRO sg13g2_nand2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2b_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 2.51 2.255 2.68 ;
        RECT 2.085 0.61 2.255 2.68 ;
        RECT 1.865 0.61 2.255 1.315 ;
        RECT 1.205 2.51 1.465 3.125 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.015 1.55 1.335 1.945 ;
    END
  END B
  PIN A_N
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.105 1.53 0.775 1.89 ;
    END
  END A_N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.715 2.935 1.975 4 ;
        RECT 0.73 2.54 0.915 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.665 -0.22 1.265 1.005 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.19 2.17 0.38 2.9 ;
      RECT 0.19 2.17 1.895 2.33 ;
      RECT 1.625 1.52 1.895 2.33 ;
      RECT 1.515 1.19 1.685 1.7 ;
      RECT 0.155 1.19 1.685 1.35 ;
      RECT 0.155 0.92 0.415 1.35 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2b_1

MACRO sg13g2_nand2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand2b_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1248 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 2.145 2.98 3.18 ;
        RECT 2.77 1 2.98 3.18 ;
        RECT 2.71 1 2.98 1.39 ;
        RECT 1.67 2.145 2.98 2.36 ;
        RECT 1.67 2.145 1.93 3.18 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 1.575 2.59 1.925 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.22 2.125 3.48 4 ;
        RECT 2.18 2.9 2.44 4 ;
        RECT 1.15 2.125 1.41 4 ;
        RECT 0.13 2.08 0.39 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 1.68 -0.22 1.94 0.855 ;
        RECT 0.13 -0.22 0.39 1.275 ;
    END
  END VSS
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.155 1.475 0.61 1.865 ;
    END
  END A_N
  OBS
    LAYER Metal1 ;
      RECT 3.2 0.53 3.48 1.2 ;
      RECT 1.155 1.035 2.45 1.2 ;
      RECT 2.18 0.53 2.45 1.2 ;
      RECT 1.155 0.5 1.415 1.2 ;
      RECT 2.18 0.53 3.48 0.76 ;
      RECT 0.64 2.08 0.9 2.88 ;
      RECT 0.805 1.015 0.965 2.34 ;
      RECT 0.805 1.585 1.47 1.845 ;
      RECT 0.64 1.015 0.965 1.275 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand2b_2

MACRO sg13g2_nand3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand3_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.95 1.57 1.325 2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.57 0.69 1.985 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.535 1.55 1.87 1.99 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1357 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 2.17 2.26 3.27 ;
        RECT 2.05 0.62 2.26 3.27 ;
        RECT 1.87 0.62 2.26 1.36 ;
        RECT 1.77 0.62 2.26 1.01 ;
        RECT 0.79 2.18 2.26 2.395 ;
        RECT 0.79 2.18 1.05 3.2 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.3 2.575 1.56 4 ;
        RECT 0.28 2.17 0.54 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.225 -0.22 0.495 0.96 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand3_1

MACRO sg13g2_nand3b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand3b_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 1.57 2.25 2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.35 1.57 1.68 1.985 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1468 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.64 2.1 3.13 3.2 ;
        RECT 2.96 0.62 3.13 3.2 ;
        RECT 2.77 0.62 3.13 1.36 ;
        RECT 2.63 0.62 3.13 1.01 ;
        RECT 1.65 2.2 3.13 2.39 ;
        RECT 1.65 2.2 1.91 3.13 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.16 2.575 2.42 4 ;
        RECT 1.14 2.17 1.4 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 1.08 -0.22 1.35 0.96 ;
    END
  END VSS
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 1.57 1.17 1.985 ;
    END
  END A_N
  OBS
    LAYER Metal1 ;
      RECT 0.44 2.235 0.86 2.86 ;
      RECT 0.44 0.88 0.61 2.86 ;
      RECT 2.43 1.54 2.78 1.87 ;
      RECT 2.43 1.2 2.59 1.87 ;
      RECT 0.44 1.2 2.59 1.37 ;
      RECT 0.44 0.88 0.71 1.37 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand3b_1

MACRO sg13g2_nand4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nand4_1 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 1.55 1.83 2 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.95 1.55 1.32 2 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.01 1.55 2.28 2 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1028 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 2.18 2.7 2.395 ;
        RECT 2.46 0.63 2.7 2.395 ;
        RECT 2.32 0.63 2.7 1.33 ;
        RECT 1.81 2.18 2.07 3.225 ;
        RECT 0.79 2.18 1.05 3.225 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.32 2.575 2.58 4 ;
        RECT 1.3 2.575 1.56 4 ;
        RECT 0.28 2.18 0.54 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 0.225 -0.22 0.495 1.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.55 0.69 2 ;
    END
  END D
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nand4_1

MACRO sg13g2_nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2_1 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.35 1.52 0.68 2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 1.52 1.54 2 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 2.235 1.54 3.125 ;
        RECT 0.87 2.235 1.54 2.435 ;
        RECT 0.87 0.605 1.135 1.35 ;
        RECT 0.87 0.605 1.04 2.435 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.4 2.24 0.66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 1.42 -0.22 1.68 1.285 ;
        RECT 0.4 -0.22 0.66 1.285 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2_1

MACRO sg13g2_nor2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.52 1.105 1.825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 1.52 2.125 1.825 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.988 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 2.055 2.6 2.36 ;
        RECT 2.345 1.075 2.6 2.36 ;
        RECT 0.81 1.075 2.6 1.315 ;
        RECT 1.78 2.055 2.13 2.64 ;
        RECT 1.83 0.59 2.085 1.315 ;
        RECT 0.81 0.59 1.065 1.315 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 0.81 2.545 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.34 -0.22 2.6 0.865 ;
        RECT 1.32 -0.22 1.58 0.865 ;
        RECT 0.3 -0.22 0.56 1.32 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.32 2.865 2.6 3.2 ;
      RECT 2.34 2.545 2.6 3.2 ;
      RECT 0.3 2.055 0.56 3.175 ;
      RECT 1.32 2.055 1.58 3.2 ;
      RECT 0.3 2.055 1.58 2.365 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2_2

MACRO sg13g2_nor2b_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2b_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.71 1.52 2.03 2 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.27 1.5 0.57 1.87 ;
    END
  END B_N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 2.235 2.03 3.125 ;
        RECT 1.36 2.235 2.03 2.435 ;
        RECT 1.36 0.605 1.625 1.35 ;
        RECT 1.36 0.605 1.53 2.435 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 0.89 2.555 1.15 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.91 -0.22 2.17 1.285 ;
        RECT 0.89 -0.22 1.15 0.87 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.25 2.08 0.51 2.88 ;
      RECT 0.25 2.08 1.15 2.26 ;
      RECT 0.89 1.05 1.15 2.26 ;
      RECT 0.25 1.05 1.15 1.31 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2b_1

MACRO sg13g2_nor2b_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor2b_2 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4784 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.17 1.54 2.96 1.825 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 0.4 0.63 0.96 ;
    END
  END B_N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9728 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.32 1.16 2.6 1.36 ;
        RECT 2.34 0.72 2.6 1.36 ;
        RECT 1.83 2 2.09 2.9 ;
        RECT 1.36 2 2.09 2.2 ;
        RECT 1.36 0.72 1.58 2.2 ;
        RECT 1.32 0.72 1.58 1.36 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 2.85 2.08 3.11 4 ;
        RECT 0.81 2.08 1.07 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.85 -0.22 3.11 1.36 ;
        RECT 1.83 -0.22 2.09 0.98 ;
        RECT 0.81 -0.22 1.07 1.42 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.32 3.08 2.6 3.26 ;
      RECT 2.34 2.08 2.6 3.26 ;
      RECT 1.32 2.475 1.58 3.26 ;
      RECT 0.27 1.16 0.53 3.04 ;
      RECT 0.27 1.705 1.18 1.865 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor2b_2

MACRO sg13g2_nor3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor3_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2457 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 1.46 0.58 2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2457 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.15 1.535 1.535 1.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2457 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.535 2.095 1.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9814 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 1.1 2.225 1.35 ;
        RECT 1.965 0.655 2.225 1.35 ;
        RECT 1.785 2.17 2.045 3.13 ;
        RECT 0.79 2.17 2.045 2.665 ;
        RECT 0.945 0.655 1.205 1.35 ;
        RECT 0.79 1.1 0.965 2.665 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 0.36 2.205 0.61 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.455 -0.22 1.715 0.845 ;
        RECT 0.36 -0.22 0.585 1.235 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor3_1

MACRO sg13g2_nor3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor3_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.485 1.575 1.295 1.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.595 1.575 2.075 1.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.82 1.575 4.165 1.9 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2692 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.31 0.72 3.57 2.765 ;
        RECT 2.29 1.6 3.57 1.86 ;
        RECT 2.29 0.72 2.55 1.86 ;
        RECT 0.76 1.175 2.55 1.375 ;
        RECT 0.76 0.72 1.02 1.375 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 1.27 2.52 1.53 4 ;
        RECT 0.25 2.08 0.51 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.325 0.22 ;
        RECT 3.82 -0.22 4.08 1.375 ;
        RECT 2.8 -0.22 3.06 1.42 ;
        RECT 1.27 -0.22 2.04 0.98 ;
        RECT 0.25 -0.22 0.51 1.375 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.78 2.945 4.08 3.205 ;
      RECT 3.82 2.08 4.08 3.205 ;
      RECT 2.8 2.08 3.06 3.205 ;
      RECT 1.78 2.52 2.04 3.205 ;
      RECT 0.76 2.125 1.02 3.16 ;
      RECT 2.29 2.125 2.55 2.765 ;
      RECT 0.76 2.125 2.55 2.34 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor3_2

MACRO sg13g2_nor4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor4_1 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 1.415 0.63 1.83 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 1.57 1.26 3.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 1.57 1.74 2.37 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 1.57 2.32 1.98 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9656 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.225 2.17 2.7 3.2 ;
        RECT 2.505 1.175 2.7 3.2 ;
        RECT 0.81 1.175 2.7 1.39 ;
        RECT 1.83 0.645 2.09 1.39 ;
        RECT 0.81 0.645 1.07 1.39 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 0.3 2.12 0.56 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.34 -0.22 2.6 0.965 ;
        RECT 1.32 -0.22 1.58 0.995 ;
        RECT 0.29 -0.22 0.56 1.23 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor4_1

MACRO sg13g2_nor4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_nor4_2 0 0 ;
  SIZE 5.76 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.485 1.575 1.295 1.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.015 1.575 2.825 1.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 1.575 3.845 1.9 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5504 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.84 0.72 5.1 2.765 ;
        RECT 0.76 1.175 5.1 1.375 ;
        RECT 3.31 0.72 3.57 1.375 ;
        RECT 2.29 0.72 2.55 1.375 ;
        RECT 0.76 0.72 1.02 1.375 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 5.76 4 ;
        RECT 1.27 2.52 1.53 4 ;
        RECT 0.25 2.08 0.51 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 5.76 0.22 ;
        RECT 5.35 -0.22 5.61 1.42 ;
        RECT 3.82 -0.22 4.59 0.98 ;
        RECT 2.8 -0.22 3.06 0.98 ;
        RECT 1.27 -0.22 2.04 0.98 ;
        RECT 0.25 -0.22 0.51 1.375 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4836 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.025 1.575 4.66 1.9 ;
    END
  END D
  OBS
    LAYER Metal1 ;
      RECT 4.33 2.945 5.61 3.205 ;
      RECT 5.35 2.08 5.61 3.205 ;
      RECT 4.33 2.125 4.59 3.205 ;
      RECT 3.31 2.125 3.57 2.765 ;
      RECT 3.31 2.125 4.59 2.305 ;
      RECT 1.78 2.945 4.08 3.205 ;
      RECT 3.82 2.505 4.08 3.205 ;
      RECT 2.8 2.08 3.06 3.205 ;
      RECT 1.78 2.52 2.04 3.205 ;
      RECT 0.76 2.125 1.02 3.16 ;
      RECT 2.29 2.125 2.55 2.765 ;
      RECT 0.76 2.125 2.55 2.34 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_nor4_2

MACRO sg13g2_o21ai_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_o21ai_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 1.43 1.55 2.06 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.77 2.64 1.93 4 ;
        RECT 0.18 2.3 0.34 4 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6772 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 2.27 1.93 2.43 ;
        RECT 1.77 0.55 1.93 2.43 ;
        RECT 1.24 2.27 1.4 3.28 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.71 -0.22 0.87 0.84 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.11 1.42 0.46 2.09 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.67 1.43 1.02 2.46 ;
    END
  END A2
  OBS
    LAYER Metal1 ;
      RECT 0.13 1.06 1.45 1.22 ;
      RECT 1.24 0.55 1.4 1.22 ;
      RECT 0.18 0.55 0.34 1.22 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_o21ai_1

MACRO sg13g2_or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or2_1 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 1.185 -0.22 1.445 1.05 ;
        RECT 0.13 -0.22 0.39 0.96 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 1.18 2.25 1.44 4 ;
        RECT 1.17 2.25 1.44 3.23 ;
    END
  END VDD
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6492 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.7 2.25 1.96 3.23 ;
        RECT 1.795 0.55 1.955 3.23 ;
        RECT 1.695 0.55 1.955 1.15 ;
    END
  END X
  PIN B
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 2.13 0.905 2.65 ;
        RECT 0.495 2.13 0.905 2.35 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.575 1.135 1.945 ;
    END
  END A
  OBS
    LAYER Metal1 ;
      RECT 0.13 2.53 0.39 3.23 ;
      RECT 0.13 1.16 0.315 3.23 ;
      RECT 1.355 1.315 1.615 1.58 ;
      RECT 0.13 1.23 1.52 1.395 ;
      RECT 0.13 1.16 0.9 1.395 ;
      RECT 0.64 0.8 0.9 1.395 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or2_1

MACRO sg13g2_or2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or2_2 0 0 ;
  SIZE 2.88 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.88 0.22 ;
        RECT 2.315 -0.22 2.575 1.2 ;
        RECT 1.185 -0.22 1.445 1.05 ;
        RECT 0.13 -0.22 0.39 0.96 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.88 4 ;
        RECT 2.315 2.205 2.575 4 ;
        RECT 1.18 2.25 1.44 4 ;
        RECT 1.17 2.25 1.44 3.23 ;
    END
  END VDD
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.837 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.7 2.25 1.96 3.23 ;
        RECT 1.795 0.55 1.955 3.23 ;
        RECT 1.695 0.55 1.955 1.15 ;
    END
  END X
  PIN B
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 2.13 0.905 2.65 ;
        RECT 0.495 2.13 0.905 2.35 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE ANALOG ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.575 1.135 1.945 ;
    END
  END A
  OBS
    LAYER Metal1 ;
      RECT 0.13 2.53 0.39 3.23 ;
      RECT 0.13 1.16 0.315 3.23 ;
      RECT 1.355 1.315 1.615 1.58 ;
      RECT 0.13 1.23 1.52 1.395 ;
      RECT 0.13 1.16 0.9 1.395 ;
      RECT 0.64 0.8 0.9 1.395 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or2_2

MACRO sg13g2_or3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or3_1 0 0 ;
  SIZE 3.36 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.74 1.505 2.07 1.935 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.505 1.56 1.935 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 1.505 0.835 1.935 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 2.04 3.05 3.2 ;
        RECT 2.89 0.605 3.05 3.2 ;
        RECT 2.76 0.605 3.05 1.305 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.36 4 ;
        RECT 1.85 2.475 2.45 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.36 0.22 ;
        RECT 2.255 -0.22 2.515 0.89 ;
        RECT 0.895 -0.22 1.155 0.89 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.385 2.12 0.645 2.995 ;
      RECT 0.385 2.12 2.515 2.295 ;
      RECT 2.345 1.115 2.515 2.295 ;
      RECT 2.345 1.52 2.71 1.85 ;
      RECT 0.385 1.115 2.515 1.325 ;
      RECT 0.385 1.11 1.965 1.325 ;
      RECT 1.445 0.675 1.965 1.325 ;
      RECT 0.385 0.765 0.645 1.325 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or3_1

MACRO sg13g2_or3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or3_2 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.74 1.505 2.07 1.935 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.505 1.56 1.935 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 1.505 0.835 1.935 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7142 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.89 1.485 3.64 1.855 ;
        RECT 2.7 2.04 3.05 3.2 ;
        RECT 2.89 0.605 3.05 3.2 ;
        RECT 2.76 0.605 3.05 1.305 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.27 2.035 3.53 4 ;
        RECT 1.85 2.475 2.45 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.285 -0.22 3.545 1.305 ;
        RECT 2.255 -0.22 2.515 0.89 ;
        RECT 0.895 -0.22 1.155 0.89 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.385 2.12 0.645 2.995 ;
      RECT 0.385 2.12 2.515 2.295 ;
      RECT 2.345 1.115 2.515 2.295 ;
      RECT 2.345 1.52 2.71 1.85 ;
      RECT 0.385 1.115 2.515 1.325 ;
      RECT 0.385 1.11 1.965 1.325 ;
      RECT 1.445 0.675 1.965 1.325 ;
      RECT 0.385 0.765 0.645 1.325 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or3_2

MACRO sg13g2_or4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or4_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 1.545 2.605 1.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.715 1.545 2.045 1.97 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.145 1.545 1.52 1.97 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 1.545 0.875 1.935 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 2.04 3.5 3.105 ;
        RECT 3.34 0.62 3.5 3.105 ;
        RECT 3.18 0.62 3.5 1.295 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.5 2.585 2.76 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.625 -0.22 2.885 1.01 ;
        RECT 1.455 -0.22 1.715 1 ;
        RECT 0.38 -0.22 0.64 1.145 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.42 2.19 0.68 3.12 ;
      RECT 0.42 2.19 2.955 2.38 ;
      RECT 2.785 1.195 2.955 2.38 ;
      RECT 2.785 1.52 3.16 1.85 ;
      RECT 2.785 1.195 2.995 1.85 ;
      RECT 0.92 1.195 2.995 1.365 ;
      RECT 2.145 0.855 2.345 1.365 ;
      RECT 0.92 0.855 1.12 1.365 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or4_1

MACRO sg13g2_or4_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_or4_2 0 0 ;
  SIZE 4.32 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.27 1.545 2.605 1.975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.715 1.545 2.045 1.97 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.145 1.545 1.52 1.97 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 1.545 0.875 1.935 ;
    END
  END D
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7681 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 2.04 3.5 3.11 ;
        RECT 3.34 0.62 3.5 3.11 ;
        RECT 3.18 0.62 3.5 1.295 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 4.32 4 ;
        RECT 3.72 2.065 3.98 4 ;
        RECT 2.5 2.585 2.76 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 4.32 0.22 ;
        RECT 3.69 -0.22 3.95 1.295 ;
        RECT 2.625 -0.22 2.885 1.01 ;
        RECT 1.455 -0.22 1.715 1 ;
        RECT 0.38 -0.22 0.64 1.145 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.42 2.19 0.68 3.12 ;
      RECT 0.42 2.19 2.955 2.38 ;
      RECT 2.785 1.195 2.955 2.38 ;
      RECT 2.785 1.52 3.16 1.85 ;
      RECT 2.785 1.195 2.995 1.85 ;
      RECT 0.92 1.195 2.995 1.365 ;
      RECT 2.145 0.855 2.345 1.365 ;
      RECT 0.92 0.855 1.12 1.365 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_or4_2

MACRO sg13g2_sdfbbp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sdfbbp_1 0 0 ;
  SIZE 16.8 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.145 0.59 16.535 3.12 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.59 2.005 14.95 3.135 ;
        RECT 14.78 0.61 14.95 3.135 ;
        RECT 14.52 0.61 14.95 1.19 ;
    END
  END Q_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.74 1.38 14.035 1.79 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4069 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.51 1.72 11.84 2 ;
        RECT 11.51 1.72 11.81 2.35 ;
        RECT 10.58 1.89 11.81 2.05 ;
        RECT 9.31 3.105 10.74 3.275 ;
        RECT 10.58 1.89 10.74 3.275 ;
        RECT 10.565 2.215 10.74 3.275 ;
        RECT 9.31 2.345 9.48 3.275 ;
        RECT 8.39 2.345 9.48 2.51 ;
        RECT 7.55 3.105 8.56 3.275 ;
        RECT 8.39 2.345 8.56 3.275 ;
        RECT 7.525 1.635 7.815 1.855 ;
        RECT 7.55 1.635 7.72 3.275 ;
    END
  END SET_B
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER Via1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal2 ;
      ANTENNAMAXAREACAR 1.167997 LAYER Metal2 ;
      ANTENNAMAXCUTCAR 0.261974 LAYER Via1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.68 1.62 2.05 2.055 ;
      LAYER Metal2 ;
        RECT 1.645 1.58 2.205 1.86 ;
      LAYER Via1 ;
        RECT 1.79 1.645 1.98 1.835 ;
    END
  END D
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2756 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 1.75 1.435 2.295 ;
    END
  END SCE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1378 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.51 1.355 0.84 2.325 ;
    END
  END SCD
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2418 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.885 1.38 4.34 1.85 ;
        RECT 3.92 1.155 4.34 1.85 ;
    END
  END CLK
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 16.8 4 ;
        RECT 15.645 2.455 15.905 4 ;
        RECT 14.055 2.885 14.315 4 ;
        RECT 12.765 2.88 13.025 4 ;
        RECT 10.925 3.055 11.57 4 ;
        RECT 8.815 2.695 9.075 4 ;
        RECT 6.915 2.34 7.175 4 ;
        RECT 4.5 2.455 4.68 4 ;
        RECT 2.92 2.855 3.18 4 ;
        RECT 0.85 2.86 1.11 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 16.8 0.22 ;
        RECT 15.675 -0.22 15.935 1.155 ;
        RECT 14.035 -0.22 14.295 1.14 ;
        RECT 11.34 -0.22 11.6 1.16 ;
        RECT 9.415 -0.22 9.59 1.175 ;
        RECT 7.01 -0.22 7.27 0.745 ;
        RECT 4.26 -0.22 4.46 0.635 ;
        RECT 2.185 -0.22 2.445 1.095 ;
        RECT 0.34 -0.22 0.6 1.055 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 15.17 1.555 15.375 3.07 ;
      RECT 15.17 1.555 15.645 1.885 ;
      RECT 15.17 0.705 15.355 3.07 ;
      RECT 11.93 2.66 12.205 3.145 ;
      RECT 11.99 2.195 12.205 3.145 ;
      RECT 10.92 2.66 12.205 2.87 ;
      RECT 10.92 2.23 11.25 2.87 ;
      RECT 11.99 2.485 14.375 2.645 ;
      RECT 14.215 1.42 14.375 2.645 ;
      RECT 11.99 2.195 12.67 2.645 ;
      RECT 12.51 0.875 12.67 2.645 ;
      RECT 14.215 1.42 14.55 1.75 ;
      RECT 12.34 0.875 12.67 1.125 ;
      RECT 13.34 1.975 13.795 2.305 ;
      RECT 13.34 0.93 13.5 2.305 ;
      RECT 12.9 1.38 13.5 1.865 ;
      RECT 13.34 0.93 13.815 1.14 ;
      RECT 12.87 0.515 13.13 1.17 ;
      RECT 11.85 0.515 12.11 1.155 ;
      RECT 11.85 0.515 13.13 0.695 ;
      RECT 9.83 2.31 10.38 2.895 ;
      RECT 10.21 0.935 10.38 2.895 ;
      RECT 12.05 1.345 12.33 1.75 ;
      RECT 10.21 1.55 11.25 1.71 ;
      RECT 11.085 1.345 11.25 1.71 ;
      RECT 10.21 0.935 10.44 1.71 ;
      RECT 11.085 1.345 12.33 1.525 ;
      RECT 9.71 1.755 10.03 2.125 ;
      RECT 9.71 1.535 9.93 2.125 ;
      RECT 9.77 0.455 9.93 2.125 ;
      RECT 10.645 0.455 10.905 1.36 ;
      RECT 9.77 0.455 10.905 0.615 ;
      RECT 7.925 2 8.16 2.905 ;
      RECT 7.925 2 9.47 2.16 ;
      RECT 9.075 1.535 9.47 2.16 ;
      RECT 6.77 0.955 6.975 1.65 ;
      RECT 9.075 0.955 9.235 2.16 ;
      RECT 6.77 0.955 9.235 1.115 ;
      RECT 8.255 0.87 8.515 1.115 ;
      RECT 8.795 0.52 9.055 0.775 ;
      RECT 7.71 0.52 8.005 0.775 ;
      RECT 7.71 0.52 9.055 0.68 ;
      RECT 6.065 2.465 6.58 2.67 ;
      RECT 6.42 0.825 6.58 2.67 ;
      RECT 6.42 1.995 7.33 2.16 ;
      RECT 7.16 1.295 7.33 2.16 ;
      RECT 8.04 1.295 8.37 1.785 ;
      RECT 7.16 1.295 8.37 1.455 ;
      RECT 5.955 0.825 6.58 0.985 ;
      RECT 5.955 0.725 6.22 0.985 ;
      RECT 5.585 2.075 5.785 2.92 ;
      RECT 1.88 2.255 2.15 2.825 ;
      RECT 1.88 2.255 2.495 2.455 ;
      RECT 2.29 1.28 2.495 2.455 ;
      RECT 5.585 2.075 6.24 2.235 ;
      RECT 6.08 1.225 6.24 2.235 ;
      RECT 1.36 1.28 2.85 1.44 ;
      RECT 2.67 0.455 2.85 1.44 ;
      RECT 5.54 1.225 6.24 1.385 ;
      RECT 1.36 0.895 1.62 1.44 ;
      RECT 5.54 0.7 5.73 1.385 ;
      RECT 3.92 0.815 5.73 0.975 ;
      RECT 5.425 0.7 5.73 0.975 ;
      RECT 3.92 0.455 4.08 0.975 ;
      RECT 2.67 0.455 4.08 0.625 ;
      RECT 4.96 2.095 5.36 3.14 ;
      RECT 5.19 1.155 5.36 3.14 ;
      RECT 5.19 1.58 5.9 1.88 ;
      RECT 4.77 1.155 5.36 1.335 ;
      RECT 3.97 2.04 4.185 3.16 ;
      RECT 3.535 2.04 4.7 2.21 ;
      RECT 4.53 1.54 4.7 2.21 ;
      RECT 3.535 0.87 3.695 2.21 ;
      RECT 4.53 1.54 5.005 1.87 ;
      RECT 3.535 0.87 3.74 1.21 ;
      RECT 3.47 2.47 3.675 3.145 ;
      RECT 2.675 2.47 3.675 2.64 ;
      RECT 2.675 2.03 3.215 2.64 ;
      RECT 3.03 0.885 3.215 2.64 ;
      RECT 1.355 3.105 2.66 3.275 ;
      RECT 2.4 2.83 2.66 3.275 ;
      RECT 0.34 2.505 0.6 3.12 ;
      RECT 1.355 2.505 1.555 3.275 ;
      RECT 0.34 2.505 1.555 2.675 ;
      RECT 8.58 1.38 8.885 1.785 ;
    LAYER Via1 ;
      RECT 13.09 1.595 13.28 1.785 ;
      RECT 8.685 1.52 8.875 1.71 ;
    LAYER Metal2 ;
      RECT 8.635 1.455 9 1.9 ;
      RECT 13.03 1.47 13.32 1.865 ;
      RECT 8.635 1.58 13.32 1.78 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sdfbbp_1

MACRO sg13g2_sighold
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_sighold 0 0 ;
  SIZE 2.4 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 2.4 4 ;
        RECT 0.57 3.17 1.925 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 2.4 0.22 ;
        RECT 0.555 -0.22 1.83 0.545 ;
    END
  END VSS
  PIN SH
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.204 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.955 2.045 2.41 ;
        RECT 0.585 1.765 2.045 2.025 ;
    END
  END SH
  OBS
    LAYER Metal1 ;
      RECT 0.175 1.325 0.405 2.41 ;
      RECT 0.175 1.325 1.245 1.585 ;
      RECT 0.175 0.955 0.395 2.41 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_sighold

MACRO sg13g2_slgcp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_slgcp_1 0 0 ;
  SIZE 8.16 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 1.865 1.525 2.37 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1807 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.38 1.51 0.785 2.18 ;
    END
  END SCE
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3978 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.585 1.575 5.89 2 ;
    END
  END CLK
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.445 2.06 7.84 3.18 ;
        RECT 7.68 0.62 7.84 3.18 ;
        RECT 7.58 0.62 7.84 1.3 ;
    END
  END GCLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 8.16 4 ;
        RECT 6.935 2.335 7.195 4 ;
        RECT 5.885 2.835 6.145 4 ;
        RECT 4.28 2.785 4.54 4 ;
        RECT 1.82 2.94 2.08 4 ;
        RECT 0.4 2.425 0.66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 8.16 0.22 ;
        RECT 7.09 -0.22 7.275 1.22 ;
        RECT 5.66 -0.22 5.92 1.275 ;
        RECT 3.99 -0.22 4.15 0.91 ;
        RECT 1.28 -0.22 1.54 0.575 ;
        RECT 0.23 -0.22 0.49 1.165 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 6.455 1.94 6.65 3.075 ;
      RECT 6.455 1.94 6.9 2.11 ;
      RECT 6.74 0.71 6.9 2.11 ;
      RECT 6.74 1.52 7.5 1.85 ;
      RECT 6.74 0.71 6.91 1.85 ;
      RECT 6.485 0.71 6.91 1.27 ;
      RECT 5.935 2.365 6.255 2.655 ;
      RECT 6.085 1.46 6.255 2.655 ;
      RECT 6.085 1.46 6.56 1.76 ;
      RECT 5.245 2.255 5.56 2.515 ;
      RECT 5.245 0.475 5.405 2.515 ;
      RECT 2.4 1.25 2.645 1.58 ;
      RECT 2.4 1.25 2.9 1.42 ;
      RECT 2.74 0.45 2.9 1.42 ;
      RECT 5.15 0.475 5.435 1.31 ;
      RECT 3.65 1.105 4.49 1.265 ;
      RECT 4.33 0.475 4.49 1.265 ;
      RECT 3.65 0.45 3.81 1.265 ;
      RECT 4.33 0.475 5.435 0.645 ;
      RECT 2.74 0.45 3.81 0.61 ;
      RECT 4.79 2 5.05 3.065 ;
      RECT 3.89 2.045 5.05 2.305 ;
      RECT 4.76 0.91 4.935 2.305 ;
      RECT 4.67 0.91 4.935 1.17 ;
      RECT 3.39 1.5 3.65 2.91 ;
      RECT 3.305 1.315 3.47 1.935 ;
      RECT 3.305 1.5 4.575 1.72 ;
      RECT 3.195 0.79 3.37 1.47 ;
      RECT 3.08 0.79 3.37 0.99 ;
      RECT 1.25 2.595 1.51 3.14 ;
      RECT 2.88 2.175 3.14 2.895 ;
      RECT 1.25 2.595 3.14 2.76 ;
      RECT 1.71 1.52 1.87 2.76 ;
      RECT 0.97 1.52 1.87 1.68 ;
      RECT 0.97 0.755 1.14 1.68 ;
      RECT 0.74 0.755 1.14 1.18 ;
      RECT 0.74 0.755 2.56 0.92 ;
      RECT 2.34 0.655 2.56 0.92 ;
      RECT 2.05 1.765 2.635 2.37 ;
      RECT 2.05 1.765 3.125 1.935 ;
      RECT 2.835 1.64 3.125 1.935 ;
      RECT 2.05 1.17 2.22 2.37 ;
      RECT 1.82 1.1 2.15 1.34 ;
    LAYER Via1 ;
      RECT 5.99 2.425 6.18 2.615 ;
      RECT 4.83 2.425 5.02 2.615 ;
    LAYER Metal2 ;
      RECT 4.76 2.42 6.255 2.62 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_slgcp_1

MACRO sg13g2_tiehi
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_tiehi 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
    END
  END VSS
  PIN L_HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3927 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 2.13 1.585 2.91 ;
    END
  END L_HI
  OBS
    LAYER Metal1 ;
      RECT 0.135 2.19 0.395 2.45 ;
      RECT 0.195 1.815 0.395 2.45 ;
      RECT 0.195 1.815 1.12 2.03 ;
      RECT 0.87 1.355 1.12 2.03 ;
      RECT 1.3 0.985 1.575 1.95 ;
      RECT 0.135 1.03 0.395 1.635 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_tiehi

MACRO sg13g2_tielo
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_tielo 0 0 ;
  SIZE 1.92 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 1.92 4 ;
        RECT 0.455 3.165 0.78 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 1.92 0.22 ;
        RECT 0.465 -0.22 0.815 0.605 ;
    END
  END VSS
  PIN L_LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2992 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.295 0.485 1.585 1.23 ;
        RECT 1.095 0.485 1.585 0.775 ;
    END
  END L_LO
  OBS
    LAYER Metal1 ;
      RECT 0.875 1.03 1.115 2.06 ;
      RECT 0.315 1.03 1.115 1.29 ;
      RECT 1.305 1.46 1.58 2.875 ;
      RECT 0.315 2.11 0.575 2.76 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_tielo

MACRO sg13g2_xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_xnor2_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7332 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.67 2.08 3.57 2.24 ;
        RECT 3.41 0.605 3.57 2.24 ;
        RECT 3.315 0.605 3.57 1.315 ;
        RECT 2.34 2.54 2.98 3.13 ;
        RECT 2.67 2.08 2.98 3.13 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4342 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.76 1.525 2.075 1.96 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4342 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.255 1.525 2.695 1.9 ;
        RECT 1.42 2.17 2.48 2.34 ;
        RECT 2.255 1.525 2.48 2.34 ;
        RECT 1.42 1.57 1.58 2.34 ;
        RECT 1.24 1.57 1.58 1.96 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 3.18 2.42 3.44 4 ;
        RECT 1.725 2.54 1.995 4 ;
        RECT 0.32 2.2 0.56 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 2.265 -0.22 2.525 0.65 ;
        RECT 0.32 -0.22 0.56 1.44 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.97 2.305 1.24 2.93 ;
      RECT 0.74 2.305 1.24 2.61 ;
      RECT 0.74 0.835 0.9 2.61 ;
      RECT 2.93 1.52 3.23 1.85 ;
      RECT 2.93 1.18 3.1 1.85 ;
      RECT 1.21 0.835 1.47 1.39 ;
      RECT 1.21 1.18 3.1 1.34 ;
      RECT 0.74 0.835 1.47 0.995 ;
      RECT 1.725 0.83 3.065 1 ;
      RECT 2.77 0.79 3.065 1 ;
      RECT 1.725 0.8 2.025 1 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_xnor2_1

MACRO sg13g2_xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sg13g2_xor2_1 0 0 ;
  SIZE 3.84 BY 3.78 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4433 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.475 1.535 2.93 1.87 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4433 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.45 0.82 1.915 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7064 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.45 2.155 3.71 3.16 ;
        RECT 3.53 1.105 3.71 3.16 ;
        RECT 2.835 1.105 3.71 1.315 ;
        RECT 2.835 0.67 3.1 1.315 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.56 3.84 4 ;
        RECT 2.43 2.895 2.69 4 ;
        RECT 0.435 2.23 0.695 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.22 3.84 0.22 ;
        RECT 3.37 -0.22 3.63 0.905 ;
        RECT 1.9 -0.22 2.16 1.34 ;
        RECT 0.285 -0.22 0.82 1.18 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 1.03 2.17 1.55 3.155 ;
      RECT 1.03 2.17 3.27 2.34 ;
      RECT 3.11 1.54 3.27 2.34 ;
      RECT 1.03 0.93 1.2 3.155 ;
      RECT 3.11 1.54 3.35 1.87 ;
      RECT 1.03 0.93 1.4 1.26 ;
      RECT 2.94 2.52 3.2 3.16 ;
      RECT 1.92 2.52 2.18 3.155 ;
      RECT 1.92 2.52 3.2 2.68 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END sg13g2_xor2_1

END LIBRARY
