*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rfcmim
C1 net1 net2 sub! rfcmim w=7u l=7u   wfeed=3u
C2 net3 net4 sub! rfcmim w=7u l=7.2u wfeed=3u
C3 net5 net6 sub! rfcmim w=7u l=7u   wfeed=5u
.ENDS
