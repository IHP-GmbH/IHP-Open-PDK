************************************************************************
* 
* Copyright 2024 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
************************************************************************


************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand3b_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand3b_1 A_N B C VDD VSS Y
*.PININFO A_N:I B:I C:I Y:O VDD:B VSS:B
MX0 net1 A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 Y net1 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 Y C VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net2 B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 net3 C VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 net1 A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 Y net1 net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

.SUBCKT sg13g2_nand3b_1_iso A_N B C VDD VSS Y
*.PININFO A_N:I B:I C:I Y:O VDD:B VSS:B
MX0 net1 A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 Y net1 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 Y C VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net2 B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 net3 C VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 net1 A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 Y net1 net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

.SUBCKT sg13g2_nand3b_1_digisub A_N B C VDD VSS Y
*.PININFO A_N:I B:I C:I Y:O VDD:B VSS:B
MX0 net1 A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 Y net1 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 Y C VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net2 B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 net3 C VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 net1 A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 Y net1 net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

