*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT pnpMPA
Q1 sub net1 net2 pnpMPA a=1.4p   p=5.4u m=1
Q2 sub net3 net4 pnpMPA a=1.5p   p=5.5u m=1
Q3 sub net5 net6 pnpMPA a=1.365p p=5.3u m=1
Q4 sub net7 net8 pnpMPA a=1.4p   p=5.4u m=3

* Extra patterns
Q_pattern_1  sub b_1  e_1  pnpMPA w=9.92u l=4.06u 
Q_pattern_2  sub b_2  e_2  pnpMPA w=1.91u l=9.91u 
Q_pattern_3  sub b_3  e_3  pnpMPA w=8.76u l=8.65u 
Q_pattern_4  sub b_4  e_4  pnpMPA w=8.38u l=4.27u 
Q_pattern_5  sub b_5  e_5  pnpMPA w=2.56u l=8.12u 
Q_pattern_6  sub b_6  e_6  pnpMPA w=1.19u l=3.38u 
Q_pattern_7  sub b_7  e_7  pnpMPA w=5.98u l=7.0u 
Q_pattern_8  sub b_8  e_8  pnpMPA w=8.88u l=8.5u 
Q_pattern_9  sub b_9  e_9  pnpMPA w=8.88u l=7.0u 
Q_pattern_10 sub b_10 e_10 pnpMPA w=5.98u l=3.38u 
Q_pattern_11 sub b_11 e_11 pnpMPA w=1.19u l=8.12u 
Q_pattern_12 sub b_12 e_12 pnpMPA w=2.56u l=4.27u 
Q_pattern_13 sub b_13 e_13 pnpMPA w=8.38u l=8.65u 
Q_pattern_14 sub b_14 e_14 pnpMPA w=8.76u l=9.91u 
Q_pattern_15 sub b_15 e_15 pnpMPA w=1.91u l=4.06u 
Q_pattern_16 sub b_16 e_16 pnpMPA w=9.92u l=8.5u 
Q_pattern_17 sub b_17 e_17 pnpMPA w=9.92u l=7.0u 
Q_pattern_18 sub b_18 e_18 pnpMPA w=1.91u l=3.38u 
Q_pattern_19 sub b_19 e_19 pnpMPA w=8.76u l=8.12u 
Q_pattern_20 sub b_20 e_20 pnpMPA w=8.38u l=8.5u 
Q_pattern_21 sub b_21 e_21 pnpMPA w=2.56u l=4.06u 
Q_pattern_22 sub b_22 e_22 pnpMPA w=1.19u l=9.91u 
Q_pattern_23 sub b_23 e_23 pnpMPA w=5.98u l=8.65u 
Q_pattern_24 sub b_24 e_24 pnpMPA w=8.88u l=4.27u 
Q_pattern_25 sub b_25 e_25 pnpMPA w=8.88u l=8.65u 
Q_pattern_26 sub b_26 e_26 pnpMPA w=5.98u l=9.91u 
Q_pattern_27 sub b_27 e_27 pnpMPA w=1.19u l=4.06u 
Q_pattern_28 sub b_28 e_28 pnpMPA w=2.56u l=8.5u 
Q_pattern_29 sub b_29 e_29 pnpMPA w=8.38u l=7.0u 
Q_pattern_30 sub b_30 e_30 pnpMPA w=8.76u l=3.38u 
Q_pattern_31 sub b_31 e_31 pnpMPA w=1.91u l=4.27u 
Q_pattern_32 sub b_32 e_32 pnpMPA w=9.92u l=8.12u 
Q_pattern_33 sub b_33 e_33 pnpMPA w=9.92u l=4.27u 
Q_pattern_34 sub b_34 e_34 pnpMPA w=1.91u l=8.65u 
Q_pattern_35 sub b_35 e_35 pnpMPA w=8.76u l=7.0u 
Q_pattern_36 sub b_36 e_36 pnpMPA w=8.38u l=4.06u 
Q_pattern_37 sub b_37 e_37 pnpMPA w=2.56u l=3.38u 
Q_pattern_38 sub b_38 e_38 pnpMPA w=1.19u l=8.5u 
Q_pattern_39 sub b_39 e_39 pnpMPA w=5.98u l=8.12u 
Q_pattern_40 sub b_40 e_40 pnpMPA w=8.88u l=9.91u 
Q_pattern_41 sub b_41 e_41 pnpMPA w=8.88u l=8.12u 
Q_pattern_42 sub b_42 e_42 pnpMPA w=5.98u l=4.06u 
Q_pattern_43 sub b_43 e_43 pnpMPA w=1.19u l=4.27u 
Q_pattern_44 sub b_44 e_44 pnpMPA w=2.56u l=7.0u 
Q_pattern_45 sub b_45 e_45 pnpMPA w=8.38u l=9.91u 
Q_pattern_46 sub b_46 e_46 pnpMPA w=8.76u l=8.5u 
Q_pattern_47 sub b_47 e_47 pnpMPA w=1.91u l=8.5u 
Q_pattern_48 sub b_48 e_48 pnpMPA w=9.92u l=3.38u 
Q_pattern_49 sub b_49 e_49 pnpMPA w=9.92u l=8.65u 
Q_pattern_50 sub b_50 e_50 pnpMPA w=1.91u l=8.12u 
Q_pattern_51 sub b_51 e_51 pnpMPA w=8.76u l=4.27u 
Q_pattern_52 sub b_52 e_52 pnpMPA w=8.38u l=3.38u 
Q_pattern_53 sub b_53 e_53 pnpMPA w=2.56u l=8.65u 
Q_pattern_54 sub b_54 e_54 pnpMPA w=1.19u l=7.0u 
Q_pattern_55 sub b_55 e_55 pnpMPA w=5.98u l=4.27u 
Q_pattern_56 sub b_56 e_56 pnpMPA w=8.88u l=4.06u 
Q_pattern_57 sub b_57 e_57 pnpMPA w=8.88u l=3.38u 
Q_pattern_58 sub b_58 e_58 pnpMPA w=5.98u l=8.5u 
Q_pattern_59 sub b_59 e_59 pnpMPA w=1.19u l=8.65u 
Q_pattern_60 sub b_60 e_60 pnpMPA w=2.56u l=9.91u 
Q_pattern_61 sub b_61 e_61 pnpMPA w=8.38u l=8.12u 
Q_pattern_62 sub b_62 e_62 pnpMPA w=8.76u l=4.06u 
Q_pattern_63 sub b_63 e_63 pnpMPA w=1.91u l=7.0u 
Q_pattern_64 sub b_64 e_64 pnpMPA w=9.92u l=9.91u 
Q_pattern_65 sub b_65 e_65 pnpMPA w=8.38u l=7.0u 
Q_pattern_66 sub b_66 e_66 pnpMPA w=1.19u l=8.5u 
.ENDS

