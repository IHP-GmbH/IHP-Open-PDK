*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT pnpMPA
Qp1 sub! net2 net3 pnpMPA a=1.4p p=5.4u m=1
Qp2 sub! net5 net6 pnpMPA a=1.5p p=5.5u m=1
Qp3 sub! net8 net9 pnpMPA a=1.365p p=5.3u m=1
Qp4 sub! net11 net12 pnpMPA a=1.4p p=5.4u m=3
.ENDS
