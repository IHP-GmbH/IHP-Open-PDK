*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT npn13G2v
QQ1 net1 net2 net3 sub! npn13G2v m=1 le=1.0u we=120.00n
QQ2 net4 net5 net6 sub! npn13G2v m=1 le=1.15u we=120.00n
QQ3 net7 net8 net9 sub! npn13G2v m=2 le=1.0u we=120.00n
.ENDS
