*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT cap_cmim
C0 PLUS1 MINUS1 $[cap_cmim] 74.620f w=6.99u l=6.99u m=1
C1 PLUS2 MINUS2 cap_cmim w=6.99u l=6.99u m=2
C2 PLUS3 MINUS3 cap_cmim w=6.99u l=6.99u m=3

* Extra patterns
C_pattern_1  plus_1  minus_1  cap_cmim w=8.1u l=18.91u 
C_pattern_2  plus_2  minus_2  cap_cmim w=16.26u l=9.81u 
C_pattern_3  plus_3  minus_3  cap_cmim w=17.93u l=18.34u 
C_pattern_4  plus_4  minus_4  cap_cmim w=17.63u l=17.92u 
C_pattern_5  plus_5  minus_5  cap_cmim w=16.97u l=11.07u 
C_pattern_6  plus_6  minus_6  cap_cmim w=15.68u l=18.27u 
C_pattern_7  plus_7  minus_7  cap_cmim w=16.88u l=11.52u 
C_pattern_8  plus_8  minus_8  cap_cmim w=9.17u l=19.85u 
C_pattern_9  plus_9  minus_9  cap_cmim w=9.17u l=11.52u 
C_pattern_10 plus_10 minus_10 cap_cmim w=16.88u l=18.27u 
C_pattern_11 plus_11 minus_11 cap_cmim w=15.68u l=11.07u 
C_pattern_12 plus_12 minus_12 cap_cmim w=16.97u l=17.92u 
C_pattern_13 plus_13 minus_13 cap_cmim w=17.63u l=18.34u 
C_pattern_14 plus_14 minus_14 cap_cmim w=17.93u l=9.81u 
C_pattern_15 plus_15 minus_15 cap_cmim w=16.26u l=18.91u 
C_pattern_16 plus_16 minus_16 cap_cmim w=8.1u l=19.85u 
C_pattern_17 plus_17 minus_17 cap_cmim w=8.1u l=11.52u 
C_pattern_18 plus_18 minus_18 cap_cmim w=16.26u l=18.27u 
C_pattern_19 plus_19 minus_19 cap_cmim w=17.93u l=11.07u 
C_pattern_20 plus_20 minus_20 cap_cmim w=17.63u l=19.85u 
C_pattern_21 plus_21 minus_21 cap_cmim w=16.97u l=18.91u 
C_pattern_22 plus_22 minus_22 cap_cmim w=15.68u l=9.81u 
C_pattern_23 plus_23 minus_23 cap_cmim w=16.88u l=18.34u 
C_pattern_24 plus_24 minus_24 cap_cmim w=9.17u l=17.92u 
C_pattern_25 plus_25 minus_25 cap_cmim w=9.17u l=18.34u 
C_pattern_26 plus_26 minus_26 cap_cmim w=16.88u l=9.81u 
C_pattern_27 plus_27 minus_27 cap_cmim w=15.68u l=18.91u 
C_pattern_28 plus_28 minus_28 cap_cmim w=16.97u l=19.85u 
C_pattern_29 plus_29 minus_29 cap_cmim w=17.63u l=11.52u 
C_pattern_30 plus_30 minus_30 cap_cmim w=17.93u l=18.27u 
C_pattern_31 plus_31 minus_31 cap_cmim w=16.26u l=17.92u 
C_pattern_32 plus_32 minus_32 cap_cmim w=8.1u l=11.07u 
C_pattern_33 plus_33 minus_33 cap_cmim w=8.1u l=17.92u 
C_pattern_34 plus_34 minus_34 cap_cmim w=16.26u l=18.34u 
C_pattern_35 plus_35 minus_35 cap_cmim w=17.93u l=11.52u 
C_pattern_36 plus_36 minus_36 cap_cmim w=17.63u l=18.91u 
C_pattern_37 plus_37 minus_37 cap_cmim w=16.97u l=18.27u 
C_pattern_38 plus_38 minus_38 cap_cmim w=15.68u l=19.85u 
C_pattern_39 plus_39 minus_39 cap_cmim w=16.88u l=11.07u 
C_pattern_40 plus_40 minus_40 cap_cmim w=9.17u l=9.81u 
C_pattern_41 plus_41 minus_41 cap_cmim w=9.17u l=11.07u 
C_pattern_42 plus_42 minus_42 cap_cmim w=16.88u l=18.91u 
C_pattern_43 plus_43 minus_43 cap_cmim w=15.68u l=17.92u 
C_pattern_44 plus_44 minus_44 cap_cmim w=16.97u l=11.52u 
C_pattern_45 plus_45 minus_45 cap_cmim w=17.63u l=9.81u 
C_pattern_46 plus_46 minus_46 cap_cmim w=17.93u l=19.85u 
C_pattern_47 plus_47 minus_47 cap_cmim w=16.26u l=19.85u 
C_pattern_48 plus_48 minus_48 cap_cmim w=8.1u l=18.27u 
C_pattern_49 plus_49 minus_49 cap_cmim w=8.1u l=18.34u 
C_pattern_50 plus_50 minus_50 cap_cmim w=16.26u l=11.07u 
C_pattern_51 plus_51 minus_51 cap_cmim w=17.93u l=17.92u 
C_pattern_52 plus_52 minus_52 cap_cmim w=17.63u l=18.27u 
C_pattern_53 plus_53 minus_53 cap_cmim w=16.97u l=18.34u 
C_pattern_54 plus_54 minus_54 cap_cmim w=15.68u l=11.52u 
C_pattern_55 plus_55 minus_55 cap_cmim w=16.88u l=17.92u 
C_pattern_56 plus_56 minus_56 cap_cmim w=9.17u l=18.91u 
C_pattern_57 plus_57 minus_57 cap_cmim w=9.17u l=18.27u 
C_pattern_58 plus_58 minus_58 cap_cmim w=16.88u l=19.85u 
C_pattern_59 plus_59 minus_59 cap_cmim w=15.68u l=18.34u 
C_pattern_60 plus_60 minus_60 cap_cmim w=16.97u l=9.81u 
C_pattern_61 plus_61 minus_61 cap_cmim w=17.63u l=11.07u 
C_pattern_62 plus_62 minus_62 cap_cmim w=17.93u l=18.91u 
C_pattern_63 plus_63 minus_63 cap_cmim w=16.26u l=11.52u 
C_pattern_64 plus_64 minus_64 cap_cmim w=8.1u l=9.81u 
C_pattern_65 plus_65 minus_65 cap_cmim w=17.63u l=11.52u 
C_pattern_66 plus_66 minus_66 cap_cmim w=15.68u l=19.85u 
.ENDS
