psp103 nch output
*
vd  d 0 dc 0.05
vg  g 0 dc 0.0
vs  s 0 dc 0.0
vb  b 0 dc 0.0
X1  d g s b sg13_lv_nmos w=1u l=0.13u mult=1

.option temp=27
.step vg 0 1.5 0.25
.dc vd 0 2.0 0.05
.print dc format=gnuplot v(d) i(vs)

.lib ../models/cornerMOSlv.lib mos_tt

.end
