*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rsil
Rs1 net1 net2 rsil m=1 l=0.5u w=0.5u
Rs2 net3 net4 rsil m=1 l=1u w=0.5u
Rs3 net5 net6 rsil m=1 l=1.2u w=0.7u
Rs4 net7 net8 rsil m=1 l=1.5u w=0.5u ps=0.2u b=1
Rs5 net9 net10 rsil m=1 l=1.7u w=0.5u ps=0.2u b=2
Rs6 net11 net12 rsil m=2 l=0.5u w=0.5u
Rs7 net13 net14 rsil m=1 l=1u w=0.5u

* Extra patterns
R_pattern_1  a_1  b_1  rsil w=5.85u l=11.25u b=3 ps=0.2u 
R_pattern_2  a_2  b_2  rsil w=1.67u l=10.81u b=6 ps=0.19u 
R_pattern_3  a_3  b_3  rsil w=4.69u l=11.80u b=4 ps=0.19u 
R_pattern_4  a_4  b_4  rsil w=5.02u l=5.84u b=4 ps=0.2u 
R_pattern_5  a_5  b_5  rsil w=0.64u l=6.94u b=2 ps=0.2u 
R_pattern_6  a_6  b_6  rsil w=4.64u l=6.62u b=4 ps=0.19u 
R_pattern_7  a_7  b_7  rsil w=3.93u l=13.27u b=8 ps=0.19u 
R_pattern_8  a_8  b_8  rsil w=5.1u l=8.13u b=9 ps=0.2u 
R_pattern_9  a_9  b_9  rsil w=5.1u l=14.44u b=4 ps=0.2u 
R_pattern_10 a_10 b_10 rsil w=3.93u l=5.91u b=2 ps=0.2u 
R_pattern_11 a_11 b_11 rsil w=4.64u l=10.94u b=4 ps=0.19u 
R_pattern_12 a_12 b_12 rsil w=0.64u l=1.46u b=4 ps=0.19u 
R_pattern_13 a_13 b_13 rsil w=5.02u l=12.13u b=6 ps=0.2u 
R_pattern_14 a_14 b_14 rsil w=4.69u l=13.83u b=3 ps=0.2u 
R_pattern_15 a_15 b_15 rsil w=1.67u l=7.07u b=9 ps=0.19u 
R_pattern_16 a_16 b_16 rsil w=5.85u l=8.88u b=8 ps=0.19u 
R_pattern_17 a_17 b_17 rsil w=1.67u l=4.70u b=2 ps=0.19u 
R_pattern_18 a_18 b_18 rsil w=5.02u l=14.36u b=4 ps=0.19u 
R_pattern_19 a_19 b_19 rsil w=4.64u l=13.78u b=8 ps=0.2u 
R_pattern_20 a_20 b_20 rsil w=5.1u l=10.50u b=4 ps=0.19u 
R_pattern_21 a_21 b_21 rsil w=5.85u l=6.67u b=6 ps=0.19u 
R_pattern_22 a_22 b_22 rsil w=4.69u l=6.67u b=9 ps=0.19u 
R_pattern_23 a_23 b_23 rsil w=0.64u l=7.75u b=3 ps=0.19u 
R_pattern_24 a_24 b_24 rsil w=3.93u l=10.23u b=4 ps=0.19u 
R_pattern_25 a_25 b_25 rsil w=1.67u l=7.97u b=4 ps=0.2u 
R_pattern_26 a_26 b_26 rsil w=3.93u l=11.04u b=4 ps=0.19u 
R_pattern_27 a_27 b_27 rsil w=0.64u l=6.04u b=4 ps=0.19u 
R_pattern_28 a_28 b_28 rsil w=4.69u l=7.72u b=4 ps=0.19u 
R_pattern_29 a_29 b_29 rsil w=5.85u l=15.19u b=2 ps=0.19u 
R_pattern_30 a_30 b_30 rsil w=5.1u l=14.24u b=2 ps=0.19u 
R_pattern_31 a_31 b_31 rsil w=4.64u l=5.46u b=9 ps=0.19u 
R_pattern_32 a_32 b_32 rsil w=5.02u l=7.00u b=3 ps=0.19u 
R_pattern_33 a_33 b_33 rsil w=5.02u l=8.05u b=8 ps=0.19u 
R_pattern_34 a_34 b_34 rsil w=4.64u l=10.04u b=6 ps=0.19u 
R_pattern_35 a_35 b_35 rsil w=5.1u l=12.21u b=8 ps=0.19u 
R_pattern_36 a_36 b_36 rsil w=5.85u l=12.15u b=9 ps=0.19u 
R_pattern_37 a_37 b_37 rsil w=4.69u l=5.51u b=2 ps=0.19u 
R_pattern_38 a_38 b_38 rsil w=0.64u l=9.98u b=9 ps=0.19u 
R_pattern_39 a_39 b_39 rsil w=3.93u l=13.07u b=9 ps=0.19u 
R_pattern_40 a_40 b_40 rsil w=1.67u l=3.65u b=4 ps=0.19u 
R_pattern_41 a_41 b_41 rsil w=1.67u l=2.49u b=3 ps=0.19u 
R_pattern_42 a_42 b_42 rsil w=3.93u l=6.96u b=6 ps=0.19u 
R_pattern_43 a_43 b_43 rsil w=0.64u l=2.62u b=6 ps=0.19u 
R_pattern_44 a_44 b_44 rsil w=4.69u l=10.09u b=8 ps=0.19u 
R_pattern_45 a_45 b_45 rsil w=5.85u l=14.99u b=4 ps=0.19u 
R_pattern_46 a_46 b_46 rsil w=5.1u l=11.40u b=3 ps=0.19u 
R_pattern_47 a_47 b_47 rsil w=4.64u l=11.75u b=2 ps=0.19u 
R_pattern_48 a_48 b_48 rsil w=5.02u l=11.32u b=4 ps=0.19u 
R_pattern_49 a_49 b_49 rsil w=5.02u l=14.16u b=4 ps=0.19u 
R_pattern_50 a_50 b_50 rsil w=4.64u l=13.98u b=3 ps=0.19u 
R_pattern_51 a_51 b_51 rsil w=5.1u l=7.08u b=4 ps=0.19u 
R_pattern_52 a_52 b_52 rsil w=5.85u l=12.96u b=4 ps=0.19u 
R_pattern_53 a_53 b_53 rsil w=4.69u l=14.03u b=4 ps=0.19u 
R_pattern_54 a_54 b_54 rsil w=0.64u l=3.67u b=4 ps=0.19u 
R_pattern_55 a_55 b_55 rsil w=3.93u l=4.75u b=4 ps=0.19u 
R_pattern_56 a_56 b_56 rsil w=1.67u l=11.01u b=6 ps=0.19u 
R_pattern_57 a_57 b_57 rsil w=5.02u l=10.42u b=2 ps=0.19u 
R_pattern_58 a_58 b_58 rsil w=1.67u l=8.78u b=9 ps=0.19u 
R_pattern_59 a_59 b_59 rsil w=4.64u l=7.67u b=4 ps=0.19u 
R_pattern_60 a_60 b_60 rsil w=1.67u l=2.49u b=8 ps=0.19u 
R_pattern_61 a_61 b_61 rsil w=3.93u l=9.33u b=3 ps=0.19u 
R_pattern_62 a_62 b_62 rsil w=0.64u l=9.78u b=8 ps=0.19u 
R_pattern_63 a_63 b_63 rsil w=4.69u l=10.99u b=6 ps=0.19u 
R_pattern_64 a_64 b_64 rsil w=5.85u l=7.83u b=4 ps=0.19u 
R_pattern_65 a_65 b_65 rsil w=5.1u l=5.92u b=6 ps=0.19u 
R_pattern_66 a_66 b_66 rsil w=5.02u l=5.84u b=9 ps=0.19u 
R_pattern_67 a_67 b_67 rsil w=1.67u l=2.49u b=4 ps=0.19u 
R_pattern_68 a_68 b_68 rsil w=5.1u l=7.08u b=8 ps=0.19u 
R_pattern_69 a_69 b_69 rsil w=5.1u l=14.24u b=4 ps=0.19u 
R_pattern_70 a_70 b_70 rsil w=5.1u l=10.50u b=4 ps=0.19u 
R_pattern_71 a_71 b_71 rsil w=5.1u l=8.13u b=4 ps=0.19u 
R_pattern_72 a_72 b_72 rsil w=5.85u l=8.88u b=3 ps=0.19u 
R_pattern_73 a_73 b_73 rsil w=4.69u l=6.67u b=4 ps=0.19u 
R_pattern_74 a_74 b_74 rsil w=0.64u l=6.94u b=8 ps=0.19u 
R_pattern_75 a_75 b_75 rsil w=3.93u l=11.04u b=4 ps=0.19u 
R_pattern_76 a_76 b_76 rsil w=3.93u l=11.04u b=2 ps=0.19u 
R_pattern_77 a_77 b_77 rsil w=3.93u l=11.04u b=4 ps=0.19u 
R_pattern_78 a_78 b_78 rsil w=4.64u l=11.75u b=4 ps=0.19u 
R_pattern_79 a_79 b_79 rsil w=5.1u l=14.44u b=4 ps=0.19u
.ENDS
