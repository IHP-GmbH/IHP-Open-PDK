*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rhigh
Rh1 net1 net2 rhigh m=1 l=0.96u w=0.5u
Rh2 net3 net4 rhigh m=1 l=1u w=0.5u
Rh3 net5 net6 rhigh m=1 l=1.2u w=0.7u
Rh4 net7 net8 rhigh m=1 l=1u w=0.5u ps=0.2u b=1
Rh5 net9 net10 rhigh m=1 l=1.2u w=0.5u ps=0.2u b=2
** Testing combiner
* res-A
R1 p_split p1 rhigh w=0.5e-6 l=30e-6 m=1 b=0
R2 p2 p_split rhigh w=0.5e-6 l=10e-6 m=1 b=0
* res-B
R3 p3 p4 rhigh w=0.5e-6 l=40e-6 m=1 b=0
* res-C with FET
R1 p5 p_intern rhigh w=0.5e-6 l=30e-6 m=1 b=0
R2 p_intern p6 rhigh w=0.5e-6 l=10e-6 m=1 b=0
M1 p_intern G S B sg13_lv_nmos w=0.15e-6 l=0.2e-6 m=1 ng=1
.ENDS
