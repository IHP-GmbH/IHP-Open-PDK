# ------------------------------------------------------
#
#		Copyright 2024 IHP PDK Authors
#
#		Licensed under the Apache License, Version 2.0 (the "License");
#		you may not use this file except in compliance with the License.
#		You may obtain a copy of the License at
#		
#		   https://www.apache.org/licenses/LICENSE-2.0
#		
#		Unless required by applicable law or agreed to in writing, software
#		distributed under the License is distributed on an "AS IS" BASIS,
#		WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
#		See the License for the specific language governing permissions and
#		limitations under the License.
#		
#		Generated on Fri Jul 19 09:01:22 2024		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_1024x8_c2_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_1024x8_c2_bm_bist 0 0 ;
  SIZE 146.88 BY 336.46 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 109.61 0 109.87 0.26 ;
    END
  END A_DIN[4]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.01 0 37.27 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 108.755 0 109.015 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 37.865 0 38.125 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 101.77 0 102.03 0.26 ;
    END
  END A_BM[4]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.85 0 45.11 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 103.145 0 103.405 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 43.475 0 43.735 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 102.28 0 102.54 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 44.34 0 44.6 0.26 ;
    END
  END A_DOUT[3]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 134.19 0 137 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.95 0 125.76 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.71 0 114.52 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 100.47 0 103.28 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 90.06 0 92.87 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 79.76 0 82.57 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.31 0 67.12 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.01 0 56.82 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 9.88 0 12.69 336.46 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 139.81 0 142.62 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.57 0 131.38 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.33 0 120.14 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.09 0 108.9 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 84.91 0 87.72 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.61 0 77.42 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 69.46 0 72.27 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.16 0 61.97 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 38.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 0 7.07 38.825 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 139.81 45.465 142.62 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.57 45.465 131.38 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 117.33 45.465 120.14 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.09 45.465 108.9 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 45.465 40.79 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 45.465 29.55 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 45.465 18.31 336.46 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.26 45.465 7.07 336.46 ;
    END
  END VDDARRAY!
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 120.85 0 121.11 0.26 ;
    END
  END A_DIN[5]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 25.77 0 26.03 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 119.995 0 120.255 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 26.625 0 26.885 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.01 0 113.27 0.26 ;
    END
  END A_BM[5]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.61 0 33.87 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 114.385 0 114.645 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 32.235 0 32.495 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 113.52 0 113.78 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 33.1 0 33.36 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 132.09 0 132.35 0.26 ;
    END
  END A_DIN[6]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 14.53 0 14.79 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 131.235 0 131.495 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 15.385 0 15.645 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.25 0 124.51 0.26 ;
    END
  END A_BM[6]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 22.37 0 22.63 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 125.625 0 125.885 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.995 0 21.255 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 124.76 0 125.02 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 21.86 0 22.12 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 143.33 0 143.59 0.26 ;
    END
  END A_DIN[7]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.838188 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 3.29 0 3.55 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 142.475 0 142.735 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6263 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.365945 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.145 0 4.405 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 135.49 0 135.75 0.26 ;
    END
  END A_BM[7]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7215 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.498382 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 11.13 0 11.39 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 136.865 0 137.125 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7605 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.055265 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 9.755 0 10.015 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 136 0 136.26 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7095 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 10.62 0 10.88 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9011 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 45.223301 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.64 0 69.9 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6967 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.184466 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 74.23 0 74.49 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.774 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 39.656958 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 69.13 0 69.39 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5696 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.618123 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 73.72 0 73.98 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 77.29 0 77.55 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 77.8 0 78.06 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 76.27 0 76.53 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6327 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 76.78 0 77.04 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1979 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.63754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 79.84 0 80.1 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9327 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.317152 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 79.33 0 79.59 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9269 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 70.245955 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.82 0 79.08 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6617 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 68.925566 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 78.31 0 78.57 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9525 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 55.436893 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.4 0 57.66 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6771 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 54.065721 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 57.91 0 58.17 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4163 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 62.724919 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 58.42 0 58.68 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1511 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.404531 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 58.93 0 59.19 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.740105 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 87.49 0 87.75 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3675 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.204381 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 88 0 88.26 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN A_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2633 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 61.963157 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.39 0 82.65 0.26 ;
    END
  END A_ADDR[9]
  PIN A_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0083 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 60.693552 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 82.9 0 83.16 0.26 ;
    END
  END A_BIST_ADDR[9]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.093851 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 67.6 0 67.86 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99505 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 20.796863 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 71.17 0 71.43 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.66 0 70.92 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0247 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.965646 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 68.11 0 68.37 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 18.532819 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 89.53 0 89.79 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9871 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 70.28015 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 10.725 LAYER Metal3 ;
      ANTENNAMAXAREACAR 3.213636 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.825655 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 70.15 0 70.41 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1639 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.953448 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 66.07 0 66.33 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1119 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 21.694548 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.7 0 72.96 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9051 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.686084 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 72.19 0 72.45 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8977 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.649241 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 66.58 0 66.84 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 146.88 336.46 ;
    LAYER Metal2 ;
      RECT 0.105 45.465 0.305 336.435 ;
      RECT 1.1 335.705 1.3 336.435 ;
      RECT 3.29 0.52 3.55 5.16 ;
      RECT 2.77 4.9 3.55 5.16 ;
      RECT 2.77 4.9 3.03 6.64 ;
      RECT 1.92 335.705 2.12 336.435 ;
      RECT 2.415 335.705 2.615 336.435 ;
      RECT 2.915 335.705 3.115 336.435 ;
      RECT 3.415 335.705 3.615 336.435 ;
      RECT 3.91 335.705 4.11 336.435 ;
      RECT 4.655 0.17 5.425 0.94 ;
      RECT 4.655 0.17 4.915 12.9 ;
      RECT 5.165 0.17 5.425 12.9 ;
      RECT 4.145 0.52 4.405 5.815 ;
      RECT 4.73 335.705 4.93 336.435 ;
      RECT 5.675 0.17 6.445 0.43 ;
      RECT 5.675 0.17 5.935 11.5 ;
      RECT 6.185 0.17 6.445 11.5 ;
      RECT 5.225 335.705 5.425 336.435 ;
      RECT 5.725 335.705 5.925 336.435 ;
      RECT 6.225 335.705 6.425 336.435 ;
      RECT 7.715 0.17 8.485 0.43 ;
      RECT 7.715 0.17 7.975 10.48 ;
      RECT 8.225 0.17 8.485 10.99 ;
      RECT 6.72 335.705 6.92 336.435 ;
      RECT 7.54 335.705 7.74 336.435 ;
      RECT 8.735 0.17 9.505 0.94 ;
      RECT 8.735 0.17 8.995 8.7 ;
      RECT 9.245 0.17 9.505 12.9 ;
      RECT 8.035 335.705 8.235 336.435 ;
      RECT 8.535 335.705 8.735 336.435 ;
      RECT 9.035 335.705 9.235 336.435 ;
      RECT 9.53 335.705 9.73 336.435 ;
      RECT 9.755 0.52 10.015 2.485 ;
      RECT 10.35 335.705 10.55 336.435 ;
      RECT 10.62 0.52 10.88 14.11 ;
      RECT 10.845 335.705 11.045 336.435 ;
      RECT 11.13 0.52 11.39 2.335 ;
      RECT 11.345 335.705 11.545 336.435 ;
      RECT 11.845 335.705 12.045 336.435 ;
      RECT 12.34 335.705 12.54 336.435 ;
      RECT 14.53 0.52 14.79 5.16 ;
      RECT 14.01 4.9 14.79 5.16 ;
      RECT 14.01 4.9 14.27 6.64 ;
      RECT 13.16 335.705 13.36 336.435 ;
      RECT 13.655 335.705 13.855 336.435 ;
      RECT 14.155 335.705 14.355 336.435 ;
      RECT 14.655 335.705 14.855 336.435 ;
      RECT 15.15 335.705 15.35 336.435 ;
      RECT 15.895 0.17 16.665 0.94 ;
      RECT 15.895 0.17 16.155 12.9 ;
      RECT 16.405 0.17 16.665 12.9 ;
      RECT 15.385 0.52 15.645 5.815 ;
      RECT 15.97 335.705 16.17 336.435 ;
      RECT 16.915 0.17 17.685 0.43 ;
      RECT 16.915 0.17 17.175 11.5 ;
      RECT 17.425 0.17 17.685 11.5 ;
      RECT 16.465 335.705 16.665 336.435 ;
      RECT 16.965 335.705 17.165 336.435 ;
      RECT 17.465 335.705 17.665 336.435 ;
      RECT 18.955 0.17 19.725 0.43 ;
      RECT 18.955 0.17 19.215 10.48 ;
      RECT 19.465 0.17 19.725 10.99 ;
      RECT 17.96 335.705 18.16 336.435 ;
      RECT 18.78 335.705 18.98 336.435 ;
      RECT 19.975 0.17 20.745 0.94 ;
      RECT 19.975 0.17 20.235 8.7 ;
      RECT 20.485 0.17 20.745 12.9 ;
      RECT 19.275 335.705 19.475 336.435 ;
      RECT 19.775 335.705 19.975 336.435 ;
      RECT 20.275 335.705 20.475 336.435 ;
      RECT 20.77 335.705 20.97 336.435 ;
      RECT 20.995 0.52 21.255 2.485 ;
      RECT 21.59 335.705 21.79 336.435 ;
      RECT 21.86 0.52 22.12 14.11 ;
      RECT 22.085 335.705 22.285 336.435 ;
      RECT 22.37 0.52 22.63 2.335 ;
      RECT 22.585 335.705 22.785 336.435 ;
      RECT 23.085 335.705 23.285 336.435 ;
      RECT 23.58 335.705 23.78 336.435 ;
      RECT 25.77 0.52 26.03 5.16 ;
      RECT 25.25 4.9 26.03 5.16 ;
      RECT 25.25 4.9 25.51 6.64 ;
      RECT 24.4 335.705 24.6 336.435 ;
      RECT 24.895 335.705 25.095 336.435 ;
      RECT 25.395 335.705 25.595 336.435 ;
      RECT 25.895 335.705 26.095 336.435 ;
      RECT 26.39 335.705 26.59 336.435 ;
      RECT 27.135 0.17 27.905 0.94 ;
      RECT 27.135 0.17 27.395 12.9 ;
      RECT 27.645 0.17 27.905 12.9 ;
      RECT 26.625 0.52 26.885 5.815 ;
      RECT 27.21 335.705 27.41 336.435 ;
      RECT 28.155 0.17 28.925 0.43 ;
      RECT 28.155 0.17 28.415 11.5 ;
      RECT 28.665 0.17 28.925 11.5 ;
      RECT 27.705 335.705 27.905 336.435 ;
      RECT 28.205 335.705 28.405 336.435 ;
      RECT 28.705 335.705 28.905 336.435 ;
      RECT 30.195 0.17 30.965 0.43 ;
      RECT 30.195 0.17 30.455 10.48 ;
      RECT 30.705 0.17 30.965 10.99 ;
      RECT 29.2 335.705 29.4 336.435 ;
      RECT 30.02 335.705 30.22 336.435 ;
      RECT 31.215 0.17 31.985 0.94 ;
      RECT 31.215 0.17 31.475 8.7 ;
      RECT 31.725 0.17 31.985 12.9 ;
      RECT 30.515 335.705 30.715 336.435 ;
      RECT 31.015 335.705 31.215 336.435 ;
      RECT 31.515 335.705 31.715 336.435 ;
      RECT 32.01 335.705 32.21 336.435 ;
      RECT 32.235 0.52 32.495 2.485 ;
      RECT 32.83 335.705 33.03 336.435 ;
      RECT 33.1 0.52 33.36 14.11 ;
      RECT 33.325 335.705 33.525 336.435 ;
      RECT 33.61 0.52 33.87 2.335 ;
      RECT 33.825 335.705 34.025 336.435 ;
      RECT 34.325 335.705 34.525 336.435 ;
      RECT 34.82 335.705 35.02 336.435 ;
      RECT 37.01 0.52 37.27 5.16 ;
      RECT 36.49 4.9 37.27 5.16 ;
      RECT 36.49 4.9 36.75 6.64 ;
      RECT 35.64 335.705 35.84 336.435 ;
      RECT 36.135 335.705 36.335 336.435 ;
      RECT 36.635 335.705 36.835 336.435 ;
      RECT 37.135 335.705 37.335 336.435 ;
      RECT 37.63 335.705 37.83 336.435 ;
      RECT 38.375 0.17 39.145 0.94 ;
      RECT 38.375 0.17 38.635 12.9 ;
      RECT 38.885 0.17 39.145 12.9 ;
      RECT 37.865 0.52 38.125 5.815 ;
      RECT 38.45 335.705 38.65 336.435 ;
      RECT 39.395 0.17 40.165 0.43 ;
      RECT 39.395 0.17 39.655 11.5 ;
      RECT 39.905 0.17 40.165 11.5 ;
      RECT 38.945 335.705 39.145 336.435 ;
      RECT 39.445 335.705 39.645 336.435 ;
      RECT 39.945 335.705 40.145 336.435 ;
      RECT 41.435 0.17 42.205 0.43 ;
      RECT 41.435 0.17 41.695 10.48 ;
      RECT 41.945 0.17 42.205 10.99 ;
      RECT 40.44 335.705 40.64 336.435 ;
      RECT 41.26 335.705 41.46 336.435 ;
      RECT 42.455 0.17 43.225 0.94 ;
      RECT 42.455 0.17 42.715 8.7 ;
      RECT 42.965 0.17 43.225 12.9 ;
      RECT 41.755 335.705 41.955 336.435 ;
      RECT 42.255 335.705 42.455 336.435 ;
      RECT 42.755 335.705 42.955 336.435 ;
      RECT 43.25 335.705 43.45 336.435 ;
      RECT 43.475 0.52 43.735 2.485 ;
      RECT 44.07 335.705 44.27 336.435 ;
      RECT 44.34 0.52 44.6 14.11 ;
      RECT 44.565 335.705 44.765 336.435 ;
      RECT 44.85 0.52 45.11 2.335 ;
      RECT 45.065 335.705 45.265 336.435 ;
      RECT 45.565 335.705 45.765 336.435 ;
      RECT 47.555 0.17 48.325 0.43 ;
      RECT 47.555 0.17 47.815 8.7 ;
      RECT 48.065 0.17 48.325 8.7 ;
      RECT 48.575 0.17 49.345 0.94 ;
      RECT 48.575 0.17 48.835 8.7 ;
      RECT 49.085 0.17 49.345 8.7 ;
      RECT 49.595 0.17 50.365 0.43 ;
      RECT 49.595 0.17 49.855 8.7 ;
      RECT 50.105 0.17 50.365 8.7 ;
      RECT 50.615 0.17 51.385 0.94 ;
      RECT 50.615 0.17 50.875 8.7 ;
      RECT 51.125 0.17 51.385 8.7 ;
      RECT 51.635 0.17 52.405 0.43 ;
      RECT 51.635 0.17 51.895 8.7 ;
      RECT 52.145 0.17 52.405 8.7 ;
      RECT 52.655 0.17 53.425 0.94 ;
      RECT 52.655 0.17 52.915 8.7 ;
      RECT 53.165 0.17 53.425 8.7 ;
      RECT 46.06 335.705 46.26 336.435 ;
      RECT 46.88 335.705 47.08 336.435 ;
      RECT 47.875 335.705 48.075 336.435 ;
      RECT 55.36 0.17 56.13 0.94 ;
      RECT 55.36 0.17 55.62 8.7 ;
      RECT 55.87 0.17 56.13 8.7 ;
      RECT 53.83 0.3 54.09 8.7 ;
      RECT 54.34 0 54.6 8.7 ;
      RECT 54.85 0 55.11 8.7 ;
      RECT 56.38 0 56.64 8.7 ;
      RECT 56.89 0 57.15 8.7 ;
      RECT 57.4 0.52 57.66 8.7 ;
      RECT 57.91 0.52 58.17 8.7 ;
      RECT 58.42 0.52 58.68 8.7 ;
      RECT 60.46 0.17 61.23 0.94 ;
      RECT 60.46 0.17 60.72 8.7 ;
      RECT 60.97 0.17 61.23 8.7 ;
      RECT 61.48 0.17 62.25 0.43 ;
      RECT 61.48 0.17 61.74 8.7 ;
      RECT 61.99 0.17 62.25 8.7 ;
      RECT 58.93 0.52 59.19 8.7 ;
      RECT 59.44 0 59.7 8.7 ;
      RECT 59.95 0 60.21 8.7 ;
      RECT 62.5 0.3 62.76 8.7 ;
      RECT 63.01 0.3 63.27 8.7 ;
      RECT 65.05 0.17 65.82 0.94 ;
      RECT 65.05 0.17 65.31 8.7 ;
      RECT 65.56 0.17 65.82 8.7 ;
      RECT 63.52 0.3 63.78 8.7 ;
      RECT 64.03 0.3 64.29 8.7 ;
      RECT 64.54 0.3 64.8 8.7 ;
      RECT 66.07 0.52 66.33 8.7 ;
      RECT 66.58 0.52 66.84 8.7 ;
      RECT 67.09 0.3 67.35 8.7 ;
      RECT 67.6 0.52 67.86 8.7 ;
      RECT 68.11 0.52 68.37 8.7 ;
      RECT 68.62 0.3 68.88 8.7 ;
      RECT 69.13 0.52 69.39 8.7 ;
      RECT 69.64 0.52 69.9 8.7 ;
      RECT 70.15 0.52 70.41 8.7 ;
      RECT 70.66 0.52 70.92 8.7 ;
      RECT 71.17 0.52 71.43 8.7 ;
      RECT 71.68 0.3 71.94 8.7 ;
      RECT 72.19 0.52 72.45 8.7 ;
      RECT 72.7 0.52 72.96 8.7 ;
      RECT 73.21 0.3 73.47 8.7 ;
      RECT 75.25 0.17 76.02 0.94 ;
      RECT 75.25 0.17 75.51 8.7 ;
      RECT 75.76 0.17 76.02 8.7 ;
      RECT 73.72 0.52 73.98 8.7 ;
      RECT 74.23 0.52 74.49 8.7 ;
      RECT 74.74 0.3 75 8.7 ;
      RECT 76.27 0.52 76.53 8.7 ;
      RECT 76.78 0.52 77.04 8.7 ;
      RECT 77.29 0.52 77.55 8.7 ;
      RECT 77.8 0.52 78.06 8.7 ;
      RECT 78.31 0.52 78.57 8.7 ;
      RECT 78.82 0.52 79.08 8.7 ;
      RECT 79.33 0.52 79.59 8.7 ;
      RECT 81.37 0.17 82.14 0.94 ;
      RECT 81.37 0.17 81.63 8.7 ;
      RECT 81.88 0.17 82.14 8.7 ;
      RECT 79.84 0.52 80.1 8.7 ;
      RECT 80.35 0 80.61 8.7 ;
      RECT 80.86 0 81.12 8.7 ;
      RECT 82.39 0.52 82.65 8.7 ;
      RECT 84.43 0.17 85.2 0.43 ;
      RECT 84.43 0.17 84.69 8.7 ;
      RECT 84.94 0.17 85.2 8.7 ;
      RECT 82.9 0.52 83.16 8.7 ;
      RECT 83.41 0.3 83.67 8.7 ;
      RECT 83.92 0.3 84.18 8.7 ;
      RECT 85.45 0.3 85.71 8.7 ;
      RECT 85.96 0.3 86.22 8.7 ;
      RECT 86.47 0.3 86.73 8.7 ;
      RECT 86.98 0.3 87.24 8.7 ;
      RECT 87.49 0.52 87.75 8.7 ;
      RECT 88 0.52 88.26 8.7 ;
      RECT 90.04 0.17 90.81 0.43 ;
      RECT 90.04 0.17 90.3 8.7 ;
      RECT 90.55 0.17 90.81 8.7 ;
      RECT 91.06 0.17 91.83 0.94 ;
      RECT 91.06 0.17 91.32 25.5 ;
      RECT 91.57 0.17 91.83 33.9 ;
      RECT 92.08 0.17 92.85 0.43 ;
      RECT 92.08 0.17 92.34 8.7 ;
      RECT 92.59 0.17 92.85 8.7 ;
      RECT 93.455 0.17 94.225 0.94 ;
      RECT 93.455 0.17 93.715 8.7 ;
      RECT 93.965 0.17 94.225 8.7 ;
      RECT 94.475 0.17 95.245 0.43 ;
      RECT 94.475 0.17 94.735 8.7 ;
      RECT 94.985 0.17 95.245 8.7 ;
      RECT 95.495 0.17 96.265 0.94 ;
      RECT 95.495 0.17 95.755 8.7 ;
      RECT 96.005 0.17 96.265 8.7 ;
      RECT 96.515 0.17 97.285 0.43 ;
      RECT 96.515 0.17 96.775 8.7 ;
      RECT 97.025 0.17 97.285 8.7 ;
      RECT 97.535 0.17 98.305 0.94 ;
      RECT 97.535 0.17 97.795 8.7 ;
      RECT 98.045 0.17 98.305 8.7 ;
      RECT 88.51 0.3 88.77 8.7 ;
      RECT 98.555 0.17 99.325 0.43 ;
      RECT 98.555 0.17 98.815 8.7 ;
      RECT 99.065 0.17 99.325 8.7 ;
      RECT 89.02 0.3 89.28 8.7 ;
      RECT 89.53 0.52 89.79 8.7 ;
      RECT 98.805 335.705 99.005 336.435 ;
      RECT 99.8 335.705 100 336.435 ;
      RECT 100.62 335.705 100.82 336.435 ;
      RECT 101.115 335.705 101.315 336.435 ;
      RECT 101.615 335.705 101.815 336.435 ;
      RECT 101.77 0.52 102.03 2.335 ;
      RECT 102.115 335.705 102.315 336.435 ;
      RECT 102.28 0.52 102.54 14.11 ;
      RECT 102.61 335.705 102.81 336.435 ;
      RECT 103.655 0.17 104.425 0.94 ;
      RECT 104.165 0.17 104.425 8.7 ;
      RECT 103.655 0.17 103.915 12.9 ;
      RECT 103.145 0.52 103.405 2.485 ;
      RECT 103.43 335.705 103.63 336.435 ;
      RECT 104.675 0.17 105.445 0.43 ;
      RECT 105.185 0.17 105.445 10.48 ;
      RECT 104.675 0.17 104.935 10.99 ;
      RECT 103.925 335.705 104.125 336.435 ;
      RECT 104.425 335.705 104.625 336.435 ;
      RECT 104.925 335.705 105.125 336.435 ;
      RECT 105.42 335.705 105.62 336.435 ;
      RECT 106.715 0.17 107.485 0.43 ;
      RECT 106.715 0.17 106.975 11.5 ;
      RECT 107.225 0.17 107.485 11.5 ;
      RECT 106.24 335.705 106.44 336.435 ;
      RECT 106.735 335.705 106.935 336.435 ;
      RECT 107.735 0.17 108.505 0.94 ;
      RECT 107.735 0.17 107.995 12.9 ;
      RECT 108.245 0.17 108.505 12.9 ;
      RECT 107.235 335.705 107.435 336.435 ;
      RECT 107.735 335.705 107.935 336.435 ;
      RECT 108.23 335.705 108.43 336.435 ;
      RECT 108.755 0.52 109.015 5.815 ;
      RECT 109.61 0.52 109.87 5.16 ;
      RECT 109.61 4.9 110.39 5.16 ;
      RECT 110.13 4.9 110.39 6.64 ;
      RECT 109.05 335.705 109.25 336.435 ;
      RECT 109.545 335.705 109.745 336.435 ;
      RECT 110.045 335.705 110.245 336.435 ;
      RECT 110.545 335.705 110.745 336.435 ;
      RECT 111.04 335.705 111.24 336.435 ;
      RECT 111.86 335.705 112.06 336.435 ;
      RECT 112.355 335.705 112.555 336.435 ;
      RECT 112.855 335.705 113.055 336.435 ;
      RECT 113.01 0.52 113.27 2.335 ;
      RECT 113.355 335.705 113.555 336.435 ;
      RECT 113.52 0.52 113.78 14.11 ;
      RECT 113.85 335.705 114.05 336.435 ;
      RECT 114.895 0.17 115.665 0.94 ;
      RECT 115.405 0.17 115.665 8.7 ;
      RECT 114.895 0.17 115.155 12.9 ;
      RECT 114.385 0.52 114.645 2.485 ;
      RECT 114.67 335.705 114.87 336.435 ;
      RECT 115.915 0.17 116.685 0.43 ;
      RECT 116.425 0.17 116.685 10.48 ;
      RECT 115.915 0.17 116.175 10.99 ;
      RECT 115.165 335.705 115.365 336.435 ;
      RECT 115.665 335.705 115.865 336.435 ;
      RECT 116.165 335.705 116.365 336.435 ;
      RECT 116.66 335.705 116.86 336.435 ;
      RECT 117.955 0.17 118.725 0.43 ;
      RECT 117.955 0.17 118.215 11.5 ;
      RECT 118.465 0.17 118.725 11.5 ;
      RECT 117.48 335.705 117.68 336.435 ;
      RECT 117.975 335.705 118.175 336.435 ;
      RECT 118.975 0.17 119.745 0.94 ;
      RECT 118.975 0.17 119.235 12.9 ;
      RECT 119.485 0.17 119.745 12.9 ;
      RECT 118.475 335.705 118.675 336.435 ;
      RECT 118.975 335.705 119.175 336.435 ;
      RECT 119.47 335.705 119.67 336.435 ;
      RECT 119.995 0.52 120.255 5.815 ;
      RECT 120.85 0.52 121.11 5.16 ;
      RECT 120.85 4.9 121.63 5.16 ;
      RECT 121.37 4.9 121.63 6.64 ;
      RECT 120.29 335.705 120.49 336.435 ;
      RECT 120.785 335.705 120.985 336.435 ;
      RECT 121.285 335.705 121.485 336.435 ;
      RECT 121.785 335.705 121.985 336.435 ;
      RECT 122.28 335.705 122.48 336.435 ;
      RECT 123.1 335.705 123.3 336.435 ;
      RECT 123.595 335.705 123.795 336.435 ;
      RECT 124.095 335.705 124.295 336.435 ;
      RECT 124.25 0.52 124.51 2.335 ;
      RECT 124.595 335.705 124.795 336.435 ;
      RECT 124.76 0.52 125.02 14.11 ;
      RECT 125.09 335.705 125.29 336.435 ;
      RECT 126.135 0.17 126.905 0.94 ;
      RECT 126.645 0.17 126.905 8.7 ;
      RECT 126.135 0.17 126.395 12.9 ;
      RECT 125.625 0.52 125.885 2.485 ;
      RECT 125.91 335.705 126.11 336.435 ;
      RECT 127.155 0.17 127.925 0.43 ;
      RECT 127.665 0.17 127.925 10.48 ;
      RECT 127.155 0.17 127.415 10.99 ;
      RECT 126.405 335.705 126.605 336.435 ;
      RECT 126.905 335.705 127.105 336.435 ;
      RECT 127.405 335.705 127.605 336.435 ;
      RECT 127.9 335.705 128.1 336.435 ;
      RECT 129.195 0.17 129.965 0.43 ;
      RECT 129.195 0.17 129.455 11.5 ;
      RECT 129.705 0.17 129.965 11.5 ;
      RECT 128.72 335.705 128.92 336.435 ;
      RECT 129.215 335.705 129.415 336.435 ;
      RECT 130.215 0.17 130.985 0.94 ;
      RECT 130.215 0.17 130.475 12.9 ;
      RECT 130.725 0.17 130.985 12.9 ;
      RECT 129.715 335.705 129.915 336.435 ;
      RECT 130.215 335.705 130.415 336.435 ;
      RECT 130.71 335.705 130.91 336.435 ;
      RECT 131.235 0.52 131.495 5.815 ;
      RECT 132.09 0.52 132.35 5.16 ;
      RECT 132.09 4.9 132.87 5.16 ;
      RECT 132.61 4.9 132.87 6.64 ;
      RECT 131.53 335.705 131.73 336.435 ;
      RECT 132.025 335.705 132.225 336.435 ;
      RECT 132.525 335.705 132.725 336.435 ;
      RECT 133.025 335.705 133.225 336.435 ;
      RECT 133.52 335.705 133.72 336.435 ;
      RECT 134.34 335.705 134.54 336.435 ;
      RECT 134.835 335.705 135.035 336.435 ;
      RECT 135.335 335.705 135.535 336.435 ;
      RECT 135.49 0.52 135.75 2.335 ;
      RECT 135.835 335.705 136.035 336.435 ;
      RECT 136 0.52 136.26 14.11 ;
      RECT 136.33 335.705 136.53 336.435 ;
      RECT 137.375 0.17 138.145 0.94 ;
      RECT 137.885 0.17 138.145 8.7 ;
      RECT 137.375 0.17 137.635 12.9 ;
      RECT 136.865 0.52 137.125 2.485 ;
      RECT 137.15 335.705 137.35 336.435 ;
      RECT 138.395 0.17 139.165 0.43 ;
      RECT 138.905 0.17 139.165 10.48 ;
      RECT 138.395 0.17 138.655 10.99 ;
      RECT 137.645 335.705 137.845 336.435 ;
      RECT 138.145 335.705 138.345 336.435 ;
      RECT 138.645 335.705 138.845 336.435 ;
      RECT 139.14 335.705 139.34 336.435 ;
      RECT 140.435 0.17 141.205 0.43 ;
      RECT 140.435 0.17 140.695 11.5 ;
      RECT 140.945 0.17 141.205 11.5 ;
      RECT 139.96 335.705 140.16 336.435 ;
      RECT 140.455 335.705 140.655 336.435 ;
      RECT 141.455 0.17 142.225 0.94 ;
      RECT 141.455 0.17 141.715 12.9 ;
      RECT 141.965 0.17 142.225 12.9 ;
      RECT 140.955 335.705 141.155 336.435 ;
      RECT 141.455 335.705 141.655 336.435 ;
      RECT 141.95 335.705 142.15 336.435 ;
      RECT 142.475 0.52 142.735 5.815 ;
      RECT 143.33 0.52 143.59 5.16 ;
      RECT 143.33 4.9 144.11 5.16 ;
      RECT 143.85 4.9 144.11 6.64 ;
      RECT 142.77 335.705 142.97 336.435 ;
      RECT 143.265 335.705 143.465 336.435 ;
      RECT 143.765 335.705 143.965 336.435 ;
      RECT 144.265 335.705 144.465 336.435 ;
      RECT 144.76 335.705 144.96 336.435 ;
      RECT 145.58 335.705 145.78 336.435 ;
      RECT 146.575 45.465 146.775 336.435 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 27.135 0.17 31.985 336.46 ;
      RECT 34.13 0 36.75 336.46 ;
      RECT 38.375 0.17 43.225 336.46 ;
      RECT 45.37 0 57.15 336.46 ;
      RECT 59.44 0.17 65.82 336.46 ;
      RECT 67.09 0.3 67.35 336.46 ;
      RECT 68.62 0.3 68.88 336.46 ;
      RECT 71.68 0.3 71.94 336.46 ;
      RECT 73.21 0.3 73.47 336.46 ;
      RECT 74.75 0.17 76.02 336.46 ;
      RECT 74.74 0.3 76.02 336.46 ;
      RECT 80.35 0.17 82.14 336.46 ;
      RECT 83.41 0.3 87.24 336.46 ;
      RECT 88.51 0.3 89.28 336.46 ;
      RECT 90.05 0 101.51 336.46 ;
      RECT 90.04 0.17 101.51 336.46 ;
      RECT 103.655 0.17 108.505 336.46 ;
      RECT 110.13 0 112.75 336.46 ;
      RECT 114.895 0.17 119.745 336.46 ;
      RECT 121.37 0 123.99 336.46 ;
      RECT 126.135 0.17 130.985 336.46 ;
      RECT 132.61 0 135.23 336.46 ;
      RECT 137.375 0.17 142.225 336.46 ;
      RECT 143.85 0 146.88 336.46 ;
      RECT 0 0.52 146.88 336.46 ;
      RECT 4.665 0 9.495 336.46 ;
      RECT 15.905 0 20.735 336.46 ;
      RECT 27.145 0 31.975 336.46 ;
      RECT 38.385 0 43.215 336.46 ;
      RECT 59.44 0 65.81 336.46 ;
      RECT 74.75 0 76.01 336.46 ;
      RECT 80.35 0 82.13 336.46 ;
      RECT 103.665 0 108.495 336.46 ;
      RECT 114.905 0 119.735 336.46 ;
      RECT 126.145 0 130.975 336.46 ;
      RECT 137.385 0 142.215 336.46 ;
      RECT 67.1 0 67.34 336.46 ;
      RECT 68.63 0 68.87 336.46 ;
      RECT 71.69 0 71.93 336.46 ;
      RECT 73.22 0 73.46 336.46 ;
      RECT 83.42 0 87.23 336.46 ;
      RECT 88.52 0 89.27 336.46 ;
      RECT 0 0 3.03 336.46 ;
      RECT 4.655 0.17 9.505 336.46 ;
      RECT 11.65 0 14.27 336.46 ;
      RECT 15.895 0.17 20.745 336.46 ;
      RECT 22.89 0 25.51 336.46 ;
    LAYER Metal3 ;
      RECT 0 0 146.88 336.46 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 0 39.085 9.62 45.205 ;
      RECT 0 0 4 336.46 ;
      RECT 7.33 0 9.62 336.46 ;
      RECT 12.95 39.085 20.86 45.205 ;
      RECT 12.95 0 15.24 336.46 ;
      RECT 18.57 0 20.86 336.46 ;
      RECT 24.19 39.085 32.1 45.205 ;
      RECT 24.19 0 26.48 336.46 ;
      RECT 29.81 0 32.1 336.46 ;
      RECT 35.43 39.085 43.34 45.205 ;
      RECT 35.43 0 37.72 336.46 ;
      RECT 41.05 0 43.34 336.46 ;
      RECT 46.67 0 53.75 336.46 ;
      RECT 57.08 0 58.9 336.46 ;
      RECT 62.23 0 64.05 336.46 ;
      RECT 67.38 0 69.2 336.46 ;
      RECT 72.53 0 74.35 336.46 ;
      RECT 77.68 0 79.5 336.46 ;
      RECT 103.54 39.085 111.45 45.205 ;
      RECT 103.54 0 105.83 336.46 ;
      RECT 109.16 0 111.45 336.46 ;
      RECT 114.78 39.085 122.69 45.205 ;
      RECT 114.78 0 117.07 336.46 ;
      RECT 120.4 0 122.69 336.46 ;
      RECT 126.02 39.085 133.93 45.205 ;
      RECT 126.02 0 128.31 336.46 ;
      RECT 131.64 0 133.93 336.46 ;
      RECT 137.26 39.085 146.88 45.205 ;
      RECT 137.26 0 139.55 336.46 ;
      RECT 142.88 0 146.88 336.46 ;
      RECT 82.83 0 84.65 336.46 ;
      RECT 87.98 0 89.8 336.46 ;
      RECT 93.13 0 100.21 336.46 ;
  END
END RM_IHPSG13_1P_1024x8_c2_bm_bist

END LIBRARY
