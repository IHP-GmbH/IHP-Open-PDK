*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT ptap1
R1 net1 sub ptap1 A=608.4f P=3.12u
R2 net2 sub ptap1 A=624.0f P=3.16u
R3 net3 sub ptap1 A=640.0f P=3.20u

* Extra patterns
R_pattern_1  a_1  sub ptap1 w=2.79u l=7.14u 
R_pattern_2  a_2  sub ptap1 w=3.42u l=7.14u 
R_pattern_3  a_3  sub ptap1 w=2.32u l=7.14u 
R_pattern_4  a_4  sub ptap1 w=8.36u l=7.14u 
R_pattern_5  a_5  sub ptap1 w=5.13u l=7.14u 
R_pattern_6  a_6  sub ptap1 w=2.4u l=7.14u 
R_pattern_7  a_7  sub ptap1 w=0.93u l=7.14u 
R_pattern_8  a_8  sub ptap1 w=3.83u l=7.14u 
R_pattern_9  a_9  sub ptap1 w=3.83u l=5.05u 
R_pattern_10 a_10 sub ptap1 w=0.93u l=5.05u 
R_pattern_11 a_11 sub ptap1 w=2.4u l=5.05u 
R_pattern_12 a_12 sub ptap1 w=5.13u l=5.05u 
R_pattern_13 a_13 sub ptap1 w=8.36u l=5.05u 
R_pattern_14 a_14 sub ptap1 w=2.32u l=5.05u 
R_pattern_15 a_15 sub ptap1 w=3.42u l=5.05u 
R_pattern_16 a_16 sub ptap1 w=2.79u l=5.05u 
R_pattern_17 a_17 sub ptap1 w=2.79u l=9.81u 
R_pattern_18 a_18 sub ptap1 w=3.42u l=9.81u 
R_pattern_19 a_19 sub ptap1 w=2.32u l=9.81u 
R_pattern_20 a_20 sub ptap1 w=8.36u l=9.81u 
R_pattern_21 a_21 sub ptap1 w=5.13u l=9.81u 
R_pattern_22 a_22 sub ptap1 w=2.4u l=9.81u 
R_pattern_23 a_23 sub ptap1 w=0.93u l=9.81u 
R_pattern_24 a_24 sub ptap1 w=3.83u l=9.81u 
R_pattern_25 a_25 sub ptap1 w=3.83u l=3.63u 
R_pattern_26 a_26 sub ptap1 w=0.93u l=3.63u 
R_pattern_27 a_27 sub ptap1 w=2.4u l=3.63u 
R_pattern_28 a_28 sub ptap1 w=5.13u l=3.63u 
R_pattern_29 a_29 sub ptap1 w=8.36u l=3.63u 
R_pattern_30 a_30 sub ptap1 w=2.32u l=3.63u 
R_pattern_31 a_31 sub ptap1 w=3.42u l=3.63u 
R_pattern_32 a_32 sub ptap1 w=2.79u l=3.63u 
R_pattern_33 a_33 sub ptap1 w=2.79u l=7.16u 
R_pattern_34 a_34 sub ptap1 w=3.42u l=7.16u 
R_pattern_35 a_35 sub ptap1 w=2.32u l=7.16u 
R_pattern_36 a_36 sub ptap1 w=8.36u l=7.16u 
R_pattern_37 a_37 sub ptap1 w=5.13u l=7.16u 
R_pattern_38 a_38 sub ptap1 w=2.4u l=7.16u 
R_pattern_39 a_39 sub ptap1 w=0.93u l=7.16u 
R_pattern_40 a_40 sub ptap1 w=3.83u l=7.16u 
R_pattern_41 a_41 sub ptap1 w=3.83u l=5.79u 
R_pattern_42 a_42 sub ptap1 w=0.93u l=5.79u 
R_pattern_43 a_43 sub ptap1 w=2.4u l=5.79u 
R_pattern_44 a_44 sub ptap1 w=5.13u l=5.79u 
R_pattern_45 a_45 sub ptap1 w=8.36u l=5.79u 
R_pattern_46 a_46 sub ptap1 w=2.32u l=5.79u 
R_pattern_47 a_47 sub ptap1 w=3.42u l=5.79u 
R_pattern_48 a_48 sub ptap1 w=2.79u l=5.79u 
R_pattern_49 a_49 sub ptap1 w=2.79u l=6.1u 
R_pattern_50 a_50 sub ptap1 w=3.42u l=6.1u 
R_pattern_51 a_51 sub ptap1 w=2.32u l=6.1u 
R_pattern_52 a_52 sub ptap1 w=8.36u l=6.1u 
R_pattern_53 a_53 sub ptap1 w=5.13u l=6.1u 
R_pattern_54 a_54 sub ptap1 w=2.4u l=6.1u 
R_pattern_55 a_55 sub ptap1 w=0.93u l=6.1u 
R_pattern_56 a_56 sub ptap1 w=3.83u l=6.1u 
R_pattern_57 a_57 sub ptap1 w=3.83u l=3.66u 
R_pattern_58 a_58 sub ptap1 w=0.93u l=3.66u 
R_pattern_59 a_59 sub ptap1 w=2.4u l=3.66u 
R_pattern_60 a_60 sub ptap1 w=5.13u l=3.66u 
R_pattern_61 a_61 sub ptap1 w=8.36u l=3.66u 
R_pattern_62 a_62 sub ptap1 w=2.32u l=3.66u 
R_pattern_63 a_63 sub ptap1 w=3.42u l=3.66u 
R_pattern_64 a_64 sub ptap1 w=2.79u l=3.66u 
.ENDS

