*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT dantenna
D1 sub net1 dantenna w=780.00n l=780.00n a=608.400f p=3.12u m=1
D2 sub net2 dantenna w=800.00n l=780.00n a=624.000f p=3.16u m=1
D3 sub net3 dantenna w=780.00n l=700.00n a=546.000f p=2.96u m=1
D4 sub net4 dantenna w=780.00n l=780.00n a=608.400f p=3.12u m=2
D5 sub net5 dantenna w=780.00n l=780.00n a=608.400f p=3.12u m=4

* Extra patterns
D_pattern_1  sub anode_1  dantenna w=9.94u l=9.73u 
D_pattern_2  sub anode_2  dantenna w=7.08u l=1.61u 
D_pattern_3  sub anode_3  dantenna w=7.11u l=5.35u 
D_pattern_4  sub anode_4  dantenna w=8.58u l=6.16u 
D_pattern_5  sub anode_5  dantenna w=9.29u l=3.88u 
D_pattern_6  sub anode_6  dantenna w=8.91u l=7.71u 
D_pattern_7  sub anode_7  dantenna w=4.93u l=6.53u 
D_pattern_8  sub anode_8  dantenna w=8.05u l=7.13u 
D_pattern_9  sub anode_9  dantenna w=8.05u l=6.53u 
D_pattern_10 sub anode_10 dantenna w=4.93u l=7.71u 
D_pattern_11 sub anode_11 dantenna w=8.91u l=3.88u 
D_pattern_12 sub anode_12 dantenna w=9.29u l=6.16u 
D_pattern_13 sub anode_13 dantenna w=8.58u l=5.35u 
D_pattern_14 sub anode_14 dantenna w=7.11u l=1.61u 
D_pattern_15 sub anode_15 dantenna w=7.08u l=9.73u 
D_pattern_16 sub anode_16 dantenna w=9.94u l=7.13u 
D_pattern_17 sub anode_17 dantenna w=9.94u l=6.53u 
D_pattern_18 sub anode_18 dantenna w=7.08u l=7.71u 
D_pattern_19 sub anode_19 dantenna w=7.11u l=3.88u 
D_pattern_20 sub anode_20 dantenna w=8.58u l=7.13u 
D_pattern_21 sub anode_21 dantenna w=9.29u l=9.73u 
D_pattern_22 sub anode_22 dantenna w=8.91u l=1.61u 
D_pattern_23 sub anode_23 dantenna w=4.93u l=5.35u 
D_pattern_24 sub anode_24 dantenna w=8.05u l=6.16u 
D_pattern_25 sub anode_25 dantenna w=8.05u l=5.35u 
D_pattern_26 sub anode_26 dantenna w=4.93u l=1.61u 
D_pattern_27 sub anode_27 dantenna w=8.91u l=9.73u 
D_pattern_28 sub anode_28 dantenna w=9.29u l=7.13u 
D_pattern_29 sub anode_29 dantenna w=8.58u l=6.53u 
D_pattern_30 sub anode_30 dantenna w=7.11u l=7.71u 
D_pattern_31 sub anode_31 dantenna w=7.08u l=6.16u 
D_pattern_32 sub anode_32 dantenna w=9.94u l=3.88u 
D_pattern_33 sub anode_33 dantenna w=9.94u l=6.16u 
D_pattern_34 sub anode_34 dantenna w=7.08u l=5.35u 
D_pattern_35 sub anode_35 dantenna w=7.11u l=6.53u 
D_pattern_36 sub anode_36 dantenna w=8.58u l=9.73u 
D_pattern_37 sub anode_37 dantenna w=9.29u l=7.71u 
D_pattern_38 sub anode_38 dantenna w=8.91u l=7.13u 
D_pattern_39 sub anode_39 dantenna w=4.93u l=3.88u 
D_pattern_40 sub anode_40 dantenna w=8.05u l=1.61u 
D_pattern_41 sub anode_41 dantenna w=8.05u l=3.88u 
D_pattern_42 sub anode_42 dantenna w=4.93u l=9.73u 
D_pattern_43 sub anode_43 dantenna w=8.91u l=6.16u 
D_pattern_44 sub anode_44 dantenna w=9.29u l=6.53u 
D_pattern_45 sub anode_45 dantenna w=8.58u l=1.61u 
D_pattern_46 sub anode_46 dantenna w=7.11u l=7.13u 
D_pattern_47 sub anode_47 dantenna w=7.08u l=7.13u 
D_pattern_48 sub anode_48 dantenna w=9.94u l=7.71u 
D_pattern_49 sub anode_49 dantenna w=9.94u l=5.35u 
D_pattern_50 sub anode_50 dantenna w=7.08u l=3.88u 
D_pattern_51 sub anode_51 dantenna w=7.11u l=6.16u 
D_pattern_52 sub anode_52 dantenna w=8.58u l=7.71u 
D_pattern_53 sub anode_53 dantenna w=9.29u l=5.35u 
D_pattern_54 sub anode_54 dantenna w=8.91u l=6.53u 
D_pattern_55 sub anode_55 dantenna w=4.93u l=6.16u 
D_pattern_56 sub anode_56 dantenna w=8.05u l=9.73u 
D_pattern_57 sub anode_57 dantenna w=8.05u l=7.71u 
D_pattern_58 sub anode_58 dantenna w=4.93u l=7.13u 
D_pattern_59 sub anode_59 dantenna w=8.91u l=5.35u 
D_pattern_60 sub anode_60 dantenna w=9.29u l=1.61u 
D_pattern_61 sub anode_61 dantenna w=8.58u l=3.88u 
D_pattern_62 sub anode_62 dantenna w=7.11u l=9.73u 
D_pattern_63 sub anode_63 dantenna w=7.08u l=6.53u 
D_pattern_64 sub anode_64 dantenna w=9.94u l=1.61u 
D_pattern_65 sub anode_65 dantenna w=8.58u l=6.53u 
D_pattern_66 sub anode_66 dantenna w=8.91u l=7.13u 
.ENDS

