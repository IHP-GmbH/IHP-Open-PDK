*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT npn13G2
Q1 C1 B1 E1 sub! npn13G2 le=900.0n we=70.00n m=1
Q2 C2 B2 E2 sub! npn13G2 le=900.0n we=70.00n m=2
Q3 C3 B3 E3 sub! npn13G2 le=900.0n we=70.00n m=4
.ENDS
