psp103 pch transfer
*
vd  d 0 dc -0.1
vg  g 0 dc 0.0
vs  s 0 dc 0.0
vb  b 0 dc 0.0
X1  d g s b sg13_lv_pmos w=1u l=0.13u mult=1
*
.option temp=27
.step vb 0 1.5 0.25
.dc vg -1.5 0.0 0.02
.print dc format=gnuplot v(g) i(vs)

.lib ../models/cornerMOSlv.lib mos_tt

.end
