*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT sg13_hv_svaricap
C1 G1 W G2 sub sg13_hv_svaricap l=0.3u w=3.74u

* Extra patterns
C_pattern_1 G1_1 W_1 G2_1 sub sg13_hv_svaricap w=7.53u l=0.36u 
C_pattern_2 G1_2 W_2 G2_2 sub sg13_hv_svaricap w=3.78u l=0.36u 
C_pattern_3 G1_3 W_3 G2_3 sub sg13_hv_svaricap w=3.78u l=0.5u 
C_pattern_4 G1_4 W_4 G2_4 sub sg13_hv_svaricap w=7.53u l=0.5u 
.ENDS
