************************************************************************
* 
* Copyright 2024 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
************************************************************************


************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_decap_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_decap_4 VDD VSS
*.PININFO VDD:B VSS:B
MX1 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
MX0 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
.ENDS

.SUBCKT sg13g2_decap_4_iso VDD VSS
*.PININFO VDD:B VSS:B
MX1 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
MX0 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
.ENDS

.SUBCKT sg13g2_decap_4_digisub VDD VSS
*.PININFO VDD:B VSS:B
MX1 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
MX0 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
.ENDS

