psp103 pch transfer
*
vd  d 0 dc -0.05
vg  g 0 dc 0.0
vs  s 0 dc 0.0
vb  b 0 dc 0.0
X1  d g s b sg13_hv_pmos w=2u l=0.5u mult=1
*
.option temp=27
.step vb 0 3 0.25
.dc vg -3 0.0 0.02
.print dc format=gnuplot v(g) i(vs)

.lib ../models/cornerMOShv.lib mos_tt

.end
