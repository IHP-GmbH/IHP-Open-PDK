*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rfcmim
C1 net1 net2 sub rfcmim w=7u l=7u   wfeed=3u
C2 net3 net4 sub rfcmim w=7.2u l=7u wfeed=3u
C3 net5 net6 sub rfcmim w=7u l=7u   wfeed=5u

* Extra patterns
C_pattern_1  plus_1  minus_1  sub rfcmim w=13.71u l=15.34u wfeed=4.13u 
C_pattern_2  plus_2  minus_2  sub rfcmim w=11.89u l=17.38u wfeed=4.13u 
C_pattern_3  plus_3  minus_3  sub rfcmim w=11.7u l=10.45u wfeed=4.13u 
C_pattern_4  plus_4  minus_4  sub rfcmim w=9.28u l=18.8u wfeed=4.13u 
C_pattern_5  plus_5  minus_5  sub rfcmim w=7.87u l=7.95u wfeed=4.13u 
C_pattern_6  plus_6  minus_6  sub rfcmim w=19.93u l=19.75u wfeed=4.13u 
C_pattern_7  plus_7  minus_7  sub rfcmim w=14.27u l=13.57u wfeed=4.13u 
C_pattern_8  plus_8  minus_8  sub rfcmim w=7.46u l=11.89u wfeed=4.13u 
C_pattern_9  plus_9  minus_9  sub rfcmim w=7.46u l=13.57u wfeed=5.87u 
C_pattern_10 plus_10 minus_10 sub rfcmim w=14.27u l=19.75u wfeed=5.87u 
C_pattern_11 plus_11 minus_11 sub rfcmim w=19.93u l=7.95u wfeed=5.87u 
C_pattern_12 plus_12 minus_12 sub rfcmim w=7.87u l=18.8u wfeed=5.87u 
C_pattern_13 plus_13 minus_13 sub rfcmim w=9.28u l=10.45u wfeed=5.87u 
C_pattern_14 plus_14 minus_14 sub rfcmim w=11.7u l=17.38u wfeed=5.87u 
C_pattern_15 plus_15 minus_15 sub rfcmim w=11.89u l=15.34u wfeed=5.87u 
C_pattern_16 plus_16 minus_16 sub rfcmim w=13.71u l=11.89u wfeed=5.87u 
C_pattern_17 plus_17 minus_17 sub rfcmim w=13.71u l=13.57u wfeed=5.61u 
C_pattern_18 plus_18 minus_18 sub rfcmim w=11.89u l=19.75u wfeed=5.61u 
C_pattern_19 plus_19 minus_19 sub rfcmim w=11.7u l=7.95u wfeed=5.61u 
C_pattern_20 plus_20 minus_20 sub rfcmim w=9.28u l=11.89u wfeed=5.61u 
C_pattern_21 plus_21 minus_21 sub rfcmim w=7.87u l=15.34u wfeed=5.61u 
C_pattern_22 plus_22 minus_22 sub rfcmim w=19.93u l=17.38u wfeed=5.61u 
C_pattern_23 plus_23 minus_23 sub rfcmim w=14.27u l=10.45u wfeed=5.61u 
C_pattern_24 plus_24 minus_24 sub rfcmim w=7.46u l=18.8u wfeed=5.61u 
C_pattern_25 plus_25 minus_25 sub rfcmim w=7.46u l=10.45u wfeed=4.89u 
C_pattern_26 plus_26 minus_26 sub rfcmim w=14.27u l=17.38u wfeed=4.89u 
C_pattern_27 plus_27 minus_27 sub rfcmim w=19.93u l=15.34u wfeed=4.89u 
C_pattern_28 plus_28 minus_28 sub rfcmim w=7.87u l=11.89u wfeed=4.89u 
C_pattern_29 plus_29 minus_29 sub rfcmim w=9.28u l=13.57u wfeed=4.89u 
C_pattern_30 plus_30 minus_30 sub rfcmim w=11.7u l=19.75u wfeed=4.89u 
C_pattern_31 plus_31 minus_31 sub rfcmim w=11.89u l=18.8u wfeed=4.89u 
C_pattern_32 plus_32 minus_32 sub rfcmim w=13.71u l=7.95u wfeed=4.89u 
C_pattern_33 plus_33 minus_33 sub rfcmim w=13.71u l=18.8u wfeed=9.9u 
C_pattern_34 plus_34 minus_34 sub rfcmim w=11.89u l=10.45u wfeed=9.9u 
C_pattern_35 plus_35 minus_35 sub rfcmim w=11.7u l=13.57u wfeed=9.9u 
C_pattern_36 plus_36 minus_36 sub rfcmim w=9.28u l=15.34u wfeed=9.9u 
C_pattern_37 plus_37 minus_37 sub rfcmim w=7.87u l=19.75u wfeed=5.12u 
C_pattern_38 plus_38 minus_38 sub rfcmim w=19.93u l=11.89u wfeed=9.9u 
C_pattern_39 plus_39 minus_39 sub rfcmim w=14.27u l=7.95u wfeed=9.9u 
C_pattern_40 plus_40 minus_40 sub rfcmim w=7.46u l=17.38u wfeed=5.12u 
C_pattern_41 plus_41 minus_41 sub rfcmim w=7.46u l=7.95u wfeed=5.69u 
C_pattern_42 plus_42 minus_42 sub rfcmim w=14.27u l=15.34u wfeed=5.12u 
C_pattern_43 plus_43 minus_43 sub rfcmim w=19.93u l=18.8u wfeed=5.69u 
C_pattern_44 plus_44 minus_44 sub rfcmim w=7.87u l=13.57u wfeed=5.69u 
C_pattern_45 plus_45 minus_45 sub rfcmim w=9.28u l=17.38u wfeed=8.47u 
C_pattern_46 plus_46 minus_46 sub rfcmim w=11.7u l=11.89u wfeed=5.69u 
C_pattern_47 plus_47 minus_47 sub rfcmim w=11.89u l=11.89u wfeed=5.12u 
C_pattern_48 plus_48 minus_48 sub rfcmim w=13.71u l=19.75u wfeed=8.47u 
C_pattern_49 plus_49 minus_49 sub rfcmim w=13.71u l=10.45u wfeed=5.69u 
C_pattern_50 plus_50 minus_50 sub rfcmim w=11.89u l=7.95u wfeed=8.47u 
C_pattern_51 plus_51 minus_51 sub rfcmim w=11.7u l=18.8u wfeed=5.12u 
C_pattern_52 plus_52 minus_52 sub rfcmim w=9.28u l=19.75u wfeed=5.69u 
C_pattern_53 plus_53 minus_53 sub rfcmim w=7.87u l=10.45u wfeed=9.9u 
C_pattern_54 plus_54 minus_54 sub rfcmim w=19.93u l=13.57u wfeed=5.12u 
C_pattern_55 plus_55 minus_55 sub rfcmim w=14.27u l=18.8u wfeed=8.47u 
C_pattern_56 plus_56 minus_56 sub rfcmim w=7.46u l=15.34u wfeed=8.47u 
C_pattern_57 plus_57 minus_57 sub rfcmim w=11.89u l=13.57u wfeed=8.47u 
C_pattern_58 plus_58 minus_58 sub rfcmim w=7.46u l=19.75u wfeed=9.9u 
C_pattern_59 plus_59 minus_59 sub rfcmim w=14.27u l=11.89u wfeed=5.69u 
C_pattern_60 plus_60 minus_60 sub rfcmim w=19.93u l=10.45u wfeed=5.12u 
C_pattern_61 plus_61 minus_61 sub rfcmim w=7.87u l=17.38u wfeed=9.9u 
C_pattern_62 plus_62 minus_62 sub rfcmim w=9.28u l=7.95u wfeed=5.12u 
C_pattern_63 plus_63 minus_63 sub rfcmim w=11.7u l=15.34u wfeed=9.9u 
C_pattern_64 plus_64 minus_64 sub rfcmim w=13.71u l=17.38u wfeed=5.69u 
C_pattern_65 plus_65 minus_65 sub rfcmim w=11.7u l=10.45u wfeed=8.47u 
C_pattern_66 plus_66 minus_66 sub rfcmim w=11.89u l=10.45u wfeed=5.69u 
C_pattern_67 plus_67 minus_67 sub rfcmim w=13.71u l=10.45u wfeed=5.12u 
C_pattern_68 plus_68 minus_68 sub rfcmim w=7.87u l=17.38u wfeed=8.47u 
C_pattern_69 plus_69 minus_69 sub rfcmim w=19.93u l=15.34u wfeed=5.12u 
C_pattern_70 plus_70 minus_70 sub rfcmim w=19.93u l=15.34u wfeed=8.47u 
C_pattern_71 plus_71 minus_71 sub rfcmim w=14.27u l=15.34u wfeed=5.69u 
C_pattern_72 plus_72 minus_72 sub rfcmim w=19.93u l=7.95u wfeed=5.12u 
C_pattern_73 plus_73 minus_73 sub rfcmim w=19.93u l=11.89u wfeed=5.69u 
C_pattern_74 plus_74 minus_74 sub rfcmim w=19.93u l=11.89u wfeed=8.47u 
C_pattern_75 plus_75 minus_75 sub rfcmim w=19.93u l=13.57u wfeed=5.69u 
C_pattern_76 plus_76 minus_76 sub rfcmim w=19.93u l=18.8u wfeed=5.69u 
.ENDS
