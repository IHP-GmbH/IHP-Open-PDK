*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT dpantenna
DD1 sub! net10 dpantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
DD2 sub! net11 dpantenna m=1 w=800.00n l=780.00n a=624.000f p=3.16u
DD3 sub! net12 dpantenna m=1 w=780.00n l=700.00n a=546.000f p=2.96u
DD4 sub! net13 dpantenna m=2 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS
