*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT inductor3
L1 net1 net2 net3 sub inductor3 w=2u s=2.1u d=25.35u nr_r=2

* Extra patterns
L_pattern_1  la__1  lc__1  lb_1  sub inductor3 w=4.49u s=9.7u d=148.305u nr_r=4
L_pattern_2  la__2  lc__2  lb_2  sub inductor3 w=8.98u s=3.74u d=151.9u nr_r=4
L_pattern_3  la__3  lc__3  lb_3  sub inductor3 w=7.54u s=5.31u d=147.605u nr_r=4
L_pattern_4  la__4  lc__4  lb_4  sub inductor3 w=4.39u s=4.96u d=103.18u nr_r=4
L_pattern_5  la__5  lc__5  lb_5  sub inductor3 w=2.9u s=8.8u d=119.235u nr_r=4
L_pattern_6  la__6  lc__6  lb_6  sub inductor3 w=4.39u s=3.74u d=52.76u nr_r=2
L_pattern_7  la__7  lc__7  lb_7  sub inductor3 w=6.96u s=3.74u d=73.955u nr_r=2
L_pattern_8  la__8  lc__8  lb_8  sub inductor3 w=8.98u s=5.31u d=97.52u nr_r=2
.ENDS
