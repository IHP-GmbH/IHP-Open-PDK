*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rhigh
Rh1 net1 net2 rhigh m=1 l=0.96u w=0.5u
Rh2 net3 net4 rhigh m=1 l=1u w=0.5u
Rh3 net5 net6 rhigh m=1 l=1.2u w=0.7u
Rh4 net7 net8 rhigh m=1 l=1u w=0.5u ps=0.2u b=1
Rh5 net9 net10 rhigh m=1 l=1.2u w=0.5u ps=0.2u b=2
** Testing combiner
* res-A
R1 p_split p1 rhigh w=0.5e-6 l=30e-6 m=1 b=0
R2 p2 p_split rhigh w=0.5e-6 l=10e-6 m=1 b=0
* res-B
R3 p3 p4 rhigh w=0.5e-6 l=40e-6 m=1 b=0
* res-C with FET
R1 p5 p_intern rhigh w=0.5e-6 l=30e-6 m=1 b=0
R2 p_intern p6 rhigh w=0.5e-6 l=10e-6 m=1 b=0
M1 p_intern G S B sg13_lv_nmos w=0.15e-6 l=0.2e-6 m=1 ng=1

* Extra patterns
R_pattern_1  a_1  b_1  rhigh w=5.85u l=5.4u b=3 ps=0.2u 
R_pattern_2  a_2  b_2  rhigh w=1.67u l=9.14u b=6 ps=0.19u 
R_pattern_3  a_3  b_3  rhigh w=4.69u l=7.11u b=4 ps=0.19u 
R_pattern_4  a_4  b_4  rhigh w=5.02u l=0.82u b=4 ps=0.2u 
R_pattern_5  a_5  b_5  rhigh w=0.64u l=6.3u b=2 ps=0.2u 
R_pattern_6  a_6  b_6  rhigh w=4.64u l=1.98u b=4 ps=0.19u 
R_pattern_7  a_7  b_7  rhigh w=3.93u l=9.34u b=8 ps=0.19u 
R_pattern_8  a_8  b_8  rhigh w=5.1u l=3.03u b=9 ps=0.2u 
R_pattern_9  a_9  b_9  rhigh w=5.1u l=9.34u b=4 ps=0.2u 
R_pattern_10 a_10 b_10 rhigh w=3.93u l=1.98u b=2 ps=0.2u 
R_pattern_11 a_11 b_11 rhigh w=4.64u l=6.3u b=4 ps=0.19u 
R_pattern_12 a_12 b_12 rhigh w=0.64u l=0.82u b=4 ps=0.19u 
R_pattern_13 a_13 b_13 rhigh w=5.02u l=7.11u b=6 ps=0.2u 
R_pattern_14 a_14 b_14 rhigh w=4.69u l=9.14u b=3 ps=0.2u 
R_pattern_15 a_15 b_15 rhigh w=1.67u l=5.4u b=9 ps=0.19u 
R_pattern_16 a_16 b_16 rhigh w=5.85u l=3.03u b=8 ps=0.19u 
R_pattern_17 a_17 b_17 rhigh w=1.67u l=3.03u b=2 ps=0.19u 
R_pattern_18 a_18 b_18 rhigh w=5.02u l=9.34u b=4 ps=0.19u 
R_pattern_19 a_19 b_19 rhigh w=4.64u l=9.14u b=8 ps=0.2u 
R_pattern_20 a_20 b_20 rhigh w=5.1u l=5.4u b=4 ps=0.19u 
R_pattern_21 a_21 b_21 rhigh w=5.85u l=0.82u b=6 ps=0.19u 
R_pattern_22 a_22 b_22 rhigh w=4.69u l=1.98u b=9 ps=0.19u 
R_pattern_23 a_23 b_23 rhigh w=0.64u l=7.11u b=3 ps=0.19u 
R_pattern_24 a_24 b_24 rhigh w=3.93u l=6.3u b=4 ps=0.19u 
R_pattern_25 a_25 b_25 rhigh w=1.67u l=6.3u b=4 ps=0.2u 
R_pattern_26 a_26 b_26 rhigh w=3.93u l=7.11u b=4 ps=0.19u 
R_pattern_27 a_27 b_27 rhigh w=0.64u l=5.4u b=4 ps=0.19u 
R_pattern_28 a_28 b_28 rhigh w=4.69u l=3.03u b=4 ps=0.19u 
R_pattern_29 a_29 b_29 rhigh w=5.85u l=9.34u b=2 ps=0.19u 
R_pattern_30 a_30 b_30 rhigh w=5.1u l=9.14u b=2 ps=0.19u 
R_pattern_31 a_31 b_31 rhigh w=4.64u l=0.82u b=9 ps=0.19u 
R_pattern_32 a_32 b_32 rhigh w=5.02u l=1.98u b=3 ps=0.19u 
R_pattern_33 a_33 b_33 rhigh w=5.02u l=3.03u b=8 ps=0.19u 
R_pattern_34 a_34 b_34 rhigh w=4.64u l=5.4u b=6 ps=0.19u 
R_pattern_35 a_35 b_35 rhigh w=5.1u l=7.11u b=8 ps=0.19u 
R_pattern_36 a_36 b_36 rhigh w=5.85u l=6.3u b=9 ps=0.19u 
R_pattern_37 a_37 b_37 rhigh w=4.69u l=0.82u b=2 ps=0.19u 
R_pattern_38 a_38 b_38 rhigh w=0.64u l=9.34u b=9 ps=0.19u 
R_pattern_39 a_39 b_39 rhigh w=3.93u l=9.14u b=9 ps=0.19u 
R_pattern_40 a_40 b_40 rhigh w=1.67u l=1.98u b=4 ps=0.19u 
R_pattern_41 a_41 b_41 rhigh w=1.67u l=0.82u b=3 ps=0.19u 
R_pattern_42 a_42 b_42 rhigh w=3.93u l=3.03u b=6 ps=0.19u 
R_pattern_43 a_43 b_43 rhigh w=0.64u l=1.98u b=6 ps=0.19u 
R_pattern_44 a_44 b_44 rhigh w=4.69u l=5.4u b=8 ps=0.19u 
R_pattern_45 a_45 b_45 rhigh w=5.85u l=9.14u b=4 ps=0.19u 
R_pattern_46 a_46 b_46 rhigh w=5.1u l=6.3u b=3 ps=0.19u 
R_pattern_47 a_47 b_47 rhigh w=4.64u l=7.11u b=2 ps=0.19u 
R_pattern_48 a_48 b_48 rhigh w=5.02u l=6.3u b=4 ps=0.19u 
R_pattern_49 a_49 b_49 rhigh w=5.02u l=9.14u b=4 ps=0.19u 
R_pattern_50 a_50 b_50 rhigh w=4.64u l=9.34u b=3 ps=0.19u 
R_pattern_51 a_51 b_51 rhigh w=5.1u l=1.98u b=4 ps=0.19u 
R_pattern_52 a_52 b_52 rhigh w=5.85u l=7.11u b=4 ps=0.19u 
R_pattern_53 a_53 b_53 rhigh w=4.69u l=9.34u b=4 ps=0.19u 
R_pattern_54 a_54 b_54 rhigh w=0.64u l=3.03u b=4 ps=0.19u 
R_pattern_55 a_55 b_55 rhigh w=3.93u l=0.82u b=4 ps=0.19u 
R_pattern_56 a_56 b_56 rhigh w=1.67u l=9.34u b=6 ps=0.19u 
R_pattern_57 a_57 b_57 rhigh w=5.02u l=5.4u b=2 ps=0.19u 
R_pattern_58 a_58 b_58 rhigh w=1.67u l=7.11u b=9 ps=0.19u 
R_pattern_59 a_59 b_59 rhigh w=4.64u l=3.03u b=4 ps=0.19u 
R_pattern_60 a_60 b_60 rhigh w=1.67u l=0.82u b=8 ps=0.19u 
R_pattern_61 a_61 b_61 rhigh w=3.93u l=5.4u b=3 ps=0.19u 
R_pattern_62 a_62 b_62 rhigh w=0.64u l=9.14u b=8 ps=0.19u 
R_pattern_63 a_63 b_63 rhigh w=4.69u l=6.3u b=6 ps=0.19u 
R_pattern_64 a_64 b_64 rhigh w=5.85u l=1.98u b=4 ps=0.19u 
R_pattern_65 a_65 b_65 rhigh w=5.1u l=0.82u b=6 ps=0.19u 
R_pattern_66 a_66 b_66 rhigh w=5.02u l=0.82u b=9 ps=0.19u 
R_pattern_67 a_67 b_67 rhigh w=1.67u l=0.82u b=4 ps=0.19u 
R_pattern_68 a_68 b_68 rhigh w=5.1u l=1.98u b=8 ps=0.19u 
R_pattern_69 a_69 b_69 rhigh w=5.1u l=9.14u b=4 ps=0.19u 
R_pattern_70 a_70 b_70 rhigh w=5.1u l=5.4u b=4 ps=0.19u 
R_pattern_71 a_71 b_71 rhigh w=5.1u l=3.03u b=4 ps=0.19u 
R_pattern_72 a_72 b_72 rhigh w=5.85u l=3.03u b=3 ps=0.19u 
R_pattern_73 a_73 b_73 rhigh w=4.69u l=1.98u b=4 ps=0.19u 
R_pattern_74 a_74 b_74 rhigh w=0.64u l=6.3u b=8 ps=0.19u 
R_pattern_75 a_75 b_75 rhigh w=3.93u l=7.11u b=4 ps=0.19u 
R_pattern_76 a_76 b_76 rhigh w=3.93u l=7.11u b=2 ps=0.19u 
R_pattern_77 a_77 b_77 rhigh w=3.93u l=7.11u b=4 ps=0.19u 
R_pattern_78 a_78 b_78 rhigh w=4.64u l=7.11u b=4 ps=0.19u 
R_pattern_79 a_79 b_79 rhigh w=5.1u l=9.34u b=4 ps=0.19u
.ENDS
