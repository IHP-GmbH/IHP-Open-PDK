*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT sg13_lv_pmos
MP1 D1 G1 S1 WELL sg13_lv_pmos w=150.00n l=130.00n ng=1 m=1
MP2 D2 G2 S2 WELL sg13_lv_pmos w=150.00n l=150.00n ng=1 m=1
MP3 D3 G3 S3 WELL sg13_lv_pmos w=200.00n l=150.00n ng=1 m=1
MP4 D4 G4 S4 WELL sg13_lv_pmos w=400.00n l=150.00n ng=2 m=1

* Extra patterns
M_pattern_37 D_37 G_37 S_37 VDD sg13_lv_pmos w=6.34u l=9.12u ng=1  
M_pattern_40 D_40 G_40 S_40 VDD sg13_lv_pmos w=5.65u l=4.99u ng=1 
M_pattern_42 D_42 G_42 S_42 VDD sg13_lv_pmos w=8.26u l=2.22u ng=1 
M_pattern_47 D_47 G_47 S_47 VDD sg13_lv_pmos w=7.15u l=0.53u ng=1 
M_pattern_51 D_51 G_51 S_51 VDD sg13_lv_pmos w=7.46u l=3.45u ng=1 
M_pattern_54 D_54 G_54 S_54 VDD sg13_lv_pmos w=9.29u l=5.38u ng=1 
M_pattern_60 D_60 G_60 S_60 VDD sg13_lv_pmos w=9.29u l=9.84u ng=1 
M_pattern_62 D_62 G_62 S_62 VDD sg13_lv_pmos w=2.74u l=4.66u ng=1 
M_pattern_67 D_67 G_67 S_67 VDD sg13_lv_pmos w=6.34u l=9.84u ng=1 
M_pattern_69 D_69 G_69 S_69 VDD sg13_lv_pmos w=9.29u l=2.22u ng=1 
M_pattern_72 D_72 G_72 S_72 VDD sg13_lv_pmos w=9.29u l=4.66u ng=1 
.ENDS
