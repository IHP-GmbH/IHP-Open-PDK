*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rfpmos
MN1 D1 G1 S1 WELL rfpmos w=1.0u l=0.72u ng=1 m=1
MN2 D2 G2 S2 WELL rfpmos w=2.0u l=0.72u ng=1 m=1
MN3 D3 G3 S3 WELL rfpmos w=1.0u l=1.0u  ng=1 m=1
MN4 D4 G4 S4 WELL rfpmos w=2.0u l=0.2u  ng=2 m=1

**** rfpmos Expected Netlist ****
M_pattern_1  D_1  G_1  S_1  VDD rfpmos w=6.93u l=2.99u ng=1 
M_pattern_2  D_2  G_2  S_2  VDD rfpmos w=3.91u l=9.48u ng=1 
M_pattern_3  D_3  G_3  S_3  VDD rfpmos w=5.66u l=5.97u ng=1 
M_pattern_4  D_4  G_4  S_4  VDD rfpmos w=6.61u l=4.57u ng=1 
M_pattern_5  D_5  G_5  S_5  VDD rfpmos w=5.7u l=8.28u ng=1 
M_pattern_6  D_6  G_6  S_6  VDD rfpmos w=9.44u l=6.89u ng=1 
M_pattern_7  D_7  G_7  S_7  VDD rfpmos w=4.34u l=9.41u ng=1 
M_pattern_8  D_8  G_8  S_8  VDD rfpmos w=2.17u l=3.22u ng=1 
M_pattern_9  D_9  G_9  S_9  VDD rfpmos w=2.17u l=9.41u ng=1 
M_pattern_10 D_10 G_10 S_10 VDD rfpmos w=4.34u l=6.89u ng=1 
M_pattern_11 D_11 G_11 S_11 VDD rfpmos w=9.44u l=8.28u ng=1 
M_pattern_12 D_12 G_12 S_12 VDD rfpmos w=5.7u l=4.57u ng=1 
M_pattern_13 D_13 G_13 S_13 VDD rfpmos w=6.61u l=5.97u ng=1 
M_pattern_14 D_14 G_14 S_14 VDD rfpmos w=5.66u l=9.48u ng=1 
M_pattern_15 D_15 G_15 S_15 VDD rfpmos w=3.91u l=2.99u ng=1 
M_pattern_16 D_16 G_16 S_16 VDD rfpmos w=6.93u l=3.22u ng=1 
.ENDS
