*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT rfnmos
MN1 D1 G1 S1 sub rfnmos w=1.0u l=0.72u ng=1 m=1
MN2 D2 G2 S2 sub rfnmos w=2.0u l=0.72u ng=1 m=1
MN3 D3 G3 S3 sub rfnmos w=1.0u l=1.0u  ng=1 m=1
MN4 D4 G4 S4 sub rfnmos w=2.0u l=0.2u  ng=2 m=1

* Extra patterns
M_pattern_37 D_37 G_37 S_37 sub rfnmos w=4.49u l=7.89u ng=1 
M_pattern_40 D_40 G_40 S_40 sub rfnmos w=6.66u l=8.06u ng=1 
M_pattern_42 D_42 G_42 S_42 sub rfnmos w=1.26u l=1.85u ng=1 
M_pattern_47 D_47 G_47 S_47 sub rfnmos w=6.58u l=5.33u ng=1 
M_pattern_51 D_51 G_51 S_51 sub rfnmos w=2.27u l=6.11u ng=1  
M_pattern_54 D_54 G_54 S_54 sub rfnmos w=8.42u l=9.74u ng=1  
M_pattern_60 D_60 G_60 S_60 sub rfnmos w=8.42u l=8.15u ng=1 
M_pattern_62 D_62 G_62 S_62 sub rfnmos w=8.83u l=6.49u ng=1 
M_pattern_67 D_67 G_67 S_67 sub rfnmos w=9.02u l=8.15u ng=1 
M_pattern_69 D_69 G_69 S_69 sub rfnmos w=8.42u l=1.85u ng=1 
M_pattern_72 D_72 G_72 S_72 sub rfnmos w=8.42u l=6.49u ng=1 
.ENDS
