*==========================================================================
* Copyright 2024 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* SPDX-License-Identifier: Apache-2.0
*==========================================================================

.SUBCKT nmos
MN1 D1 G1 S1 B sg13_lv_nmos m=1 w=150.00n l=130.00n ng=1
MN2 D2 G2 S2 B sg13_lv_nmos m=1 w=200.00n l=130.00n ng=1
MN3 D3 G3 S3 B sg13_lv_nmos m=1 w=200.00n l=150.00n ng=1
MN4 D4 G4 S4 B sg13_lv_nmos m=1 w=300.00n l=150.00n ng=2
.ENDS
